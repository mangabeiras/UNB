CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 300 100 9
0 66 421 409
7 5.000 V
7 5.000 V
3 GND
5000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 421 409
9961490 0
0
0
0
0
0
0
15
5 SAVE-
218 348 182 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
26 *Combine
*TRAN -14m 15.6m
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 71 167 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
26 *Combine
*TRAN -14m 15.6m
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
7 Ground~
168 91 210 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 348 235 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
11 Signal Gen~
195 43 172 0 19 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1176256512 0 1065353216
20
1 10000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 320 0
5 -1/1V
-17 -28 18 -20
2 V1
-7 -38 7 -30
0
0
37 %D %1 %2 DC 0 SIN(0 1 10k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
2 +V
167 207 293 0 1 3
0 8
0
0 0 53600 -19276
4 -12V
7 -7 35 1
2 V2
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
2 +V
167 209 47 0 1 3
0 9
0
0 0 53600 0
4 +12V
9 -2 37 6
2 V3
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
12 PNP Trans:C~
219 240 221 0 3 7
0 8 5 6
12 PNP Trans:C~
0 0 320 692
7 2N2905A
16 -4 65 4
2 Q1
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
4 TO-5
7

0 3 2 1 3 2 1 -33686019
113 0 0 0 1 1 0 0
1 Q
3747 0 0
0
0
12 NPN Trans:C~
219 240 114 0 3 7
0 9 7 6
12 NPN Trans:C~
0 0 320 0
7 2N2219A
16 -4 65 4
2 Q2
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
4 TO-5
7

0 3 2 1 3 2 1 -33686019
81 0 0 0 1 1 0 0
1 Q
3549 0 0
0
0
10 Capacitor~
219 113 167 0 2 5
0 4 3
10 Capacitor~
0 0 320 0
6 1.26uF
-22 -18 20 -10
2 C1
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
7931 0 0
0
0
9 Resistor~
219 152 88 0 4 5
0 7 9 0 1
9 Resistor~
0 0 352 90
3 16k
7 -5 28 3
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 152 140 0 2 5
0 3 7
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 152 194 0 2 5
0 5 3
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 152 248 0 3 5
0 8 5 1
9 Resistor~
0 0 352 90
3 16k
7 -5 28 3
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 348 197 0 3 5
0 2 6 -1
9 Resistor~
0 0 352 90
2 50
8 -5 22 3
2 R5
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
7668 0 0
0
0
15
2 0 3 0 0 4224 0 10 0 0 12 2
122 167
152 167
1 1 4 0 0 4224 0 5 10 0 0 2
74 167
104 167
2 0 5 0 0 4224 0 8 0 0 11 2
222 221
152 221
1 1 2 0 0 4096 0 15 4 0 0 2
348 215
348 229
2 0 6 0 0 8320 0 15 0 0 7 3
348 179
348 166
245 166
2 0 7 0 0 4224 0 9 0 0 13 2
222 114
152 114
3 3 6 0 0 0 0 9 8 0 0 2
245 132
245 203
1 2 2 0 0 4224 0 3 5 0 0 3
91 204
91 177
74 177
1 0 8 0 0 4096 0 6 0 0 10 2
207 278
207 270
1 1 8 0 0 8320 0 14 8 0 0 4
152 266
152 270
245 270
245 239
1 2 5 0 0 0 0 13 14 0 0 2
152 212
152 230
1 2 3 0 0 0 0 12 13 0 0 2
152 158
152 176
1 2 7 0 0 0 0 11 12 0 0 2
152 106
152 122
1 0 9 0 0 4096 0 7 0 0 15 2
209 56
209 65
2 1 9 0 0 8320 0 11 9 0 0 4
152 70
152 65
245 65
245 96
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
200 0 1 1e+006
0 0.001 2.5e-006 2.5e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2740 8550976 100 100 0 0
98 66 608 126
0 259 640 452
608 66
98 66
608 66
608 126
0 0
4.85009e-315 0 5.02117e-315 1.56312e-314 4.85009e-315 4.85009e-315
12409 0
4 0.0003 5
2
348 179
0 6 0 0 1	0 5 0 0
74 167
0 4 0 0 1	0 2 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
