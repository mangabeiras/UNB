CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
0 66 640 259
144179216 0
0
0
0
0
0
0
8
5 SAVE-
218 114 29 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
18 *DC 0.000 250.0m 0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
4 SAVE
8953 0 0
0
0
9 I Source~
198 56 92 0 2 5
0 2 3
0
0 0 16992 90
5 100mA
12 -2 47 6
3 Ibb
-11 -20 10 -12
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 0 0 0 0
2 Is
4441 0 0
0
0
9 V Source~
197 225 70 0 2 5
0 5 2
0
0 0 16992 0
3 10V
12 -2 33 6
3 Vce
13 -5 34 3
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
3618 0 0
0
0
9 V Source~
197 113 46 0 2 5
0 5 4
0
0 0 16736 0
2 0V
15 -2 29 6
3 Vs1
12 -12 33 -4
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
6153 0 0
0
0
7 Ground~
168 225 125 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 24 120 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 113 127 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
12 NPN Trans:C~
219 108 92 0 3 7
0 4 3 2
12 NPN Trans:C~
0 0 320 0
6 2N3904
20 -4 62 4
2 Q1
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 -1 261 0 1 1 0 0
1 Q
3747 0 0
0
0
6
1 1 2 0 0 4096 0 6 2 0 0 3
24 114
24 92
35 92
2 2 3 0 0 4224 0 8 2 0 0 2
90 92
77 92
3 1 2 0 0 0 0 8 7 0 0 2
113 110
113 121
2 1 4 0 0 4224 0 4 8 0 0 2
113 67
113 74
1 1 5 0 0 8320 0 3 4 0 0 4
225 49
225 6
113 6
113 25
2 1 2 0 0 4224 0 3 5 0 0 2
225 91
225 119
0
0
4 0 0
0
0
3 Vce
0 4 0.02
3 Ibb
0.001 0.01 0.002
3 0 1 4
0 2e-006 1e-008 1e-008 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
1212 2259520 100 100 0 0
98 66 608 126
0 259 640 452
608 66
98 66
608 66
608 126
0 0
5.34602e-315 0 4.99564e-315 0 5.34602e-315 4.99564e-315
12409 0
4 1 0.1
1
113 28
0 5 0 0 1	4 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
