CircuitMaker Text
5.6
Probes: 2
vin
Transient Analysis
0 269 138 65280
vout
Transient Analysis
1 425 138 65535
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
231 152 911 669
7 5.000 V
7 5.000 V
3 GND
192 10
24 100 1 1 0
20 Package,Description,
64 D:\Program Files\Protel Technology\CircuitMaker 2000 Pro\BOM.DAT
0 7
2 4 0.500000 0.500000
231 411 911 669
9961472 0
0
0
0
0
0
0
9
7 Ground~
168 327 284 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 15449516
0 0 0 0 1 0 0 0
0
9187 0 0
2
36626.6 0
0
11 Signal Gen~
195 89 130 0 19 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1114636288 1094713344 1045220557
20
1 60 12 0.2 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 49488 0
10 11.8/12.2V
-34 -29 36 -21
2 V1
-7 -38 7 -30
0
0
40 %D %1 %2 DC 0 SIN(12 200m 60 0 0) AC 1 0
0
0
0
5

0 1 2 1 2 94
86 0 0 0 1 0 0 0
1 V
6114 0 0
2
36626.6 1
0
12 NPN Trans:C~
219 329 144 0 3 64
0 4 9 3
12 NPN Trans:C~
0 0 1872 90
7 2N2222A
-26 -28 23 -20
2 Q1
-9 -40 5 -32
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 1 2 3 1 2 3 22
81 0 0 0 1 0 0 0
1 Q
7399 0 0
2
36626.6 2
0
10 Polar Cap~
219 366 205 0 2 64
0 3 2
10 Polar Cap~
0 0 1872 26894
5 100uF
13 -3 48 5
2 C1
23 -13 37 -5
0
0
11 %D %1 %2 %V
0
0
7 RB.2/.4
5

0 1 2 1 2 15490724
67 0 0 0 1 0 0 0
1 C
3374 0 0
2
36626.6 3
0
12 Zener Diode~
219 327 231 0 2 64
0 2 9
12 Zener Diode~
0 0 1872 90
6 1N4736
-57 0 -15 8
2 D1
-43 -10 -29 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 28846756
100 0 0 0 1 0 0 0
1 D
6973 0 0
2
36626.6 4
0
5 SIP2~
219 477 141 0 2 64
0 3 2
5 SIP2~
0 0 3952 0
6 Output
-22 -21 20 -13
2 J2
-8 -29 6 -21
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 15481944
0 0 0 0 1 1 0 0
1 J
5327 0 0
2
36626.6 5
0
5 SIP2~
219 208 141 0 2 64
0 4 2
5 SIP2~
0 0 3952 512
5 Input
-19 -21 16 -13
2 J1
-11 -29 3 -21
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 15514728
0 0 0 0 1 1 0 0
1 J
4244 0 0
2
36626.6 6
0
9 Resistor~
219 257 178 0 2 64
0 9 4
9 Resistor~
0 0 1904 90
3 680
7 5 28 13
2 R1
9 -5 23 3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 122
82 0 0 0 1 0 0 0
1 R
9590 0 0
2
36626.6 7
0
9 Resistor~
219 530 137 0 3 64
0 2 3 -1
9 Resistor~
0 0 49520 90
3 100
9 -5 30 3
2 RL
12 -15 26 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 15514200
82 0 0 0 1 0 0 0
1 R
5112 0 0
2
36626.6 8
0
18
0 0 5 0 0 8320 0 0 0 0 0 4
184 90
184 69
500 69
500 86
0 0 6 0 0 4224 0 0 0 0 0 2
500 177
500 101
0 0 7 0 0 8320 0 0 0 0 0 4
183 175
183 299
500 299
500 197
0 0 8 0 0 4224 0 0 0 0 0 2
184 101
184 160
0 1 2 0 0 8192 0 0 9 9 0 4
450 146
450 186
530 186
530 155
0 2 3 0 0 8192 0 0 9 17 0 4
450 137
450 93
530 93
530 119
2 0 2 0 0 0 0 2 0 0 10 5
120 135
148 135
148 166
227 166
227 146
1 0 4 0 0 12288 0 2 0 0 18 5
120 125
148 125
148 95
227 95
227 137
2 0 2 0 0 8320 0 6 0 0 13 4
465 146
438 146
438 258
365 258
2 0 2 0 0 0 0 7 0 0 14 4
214 146
239 146
239 258
327 258
1 0 9 0 0 8320 0 8 0 0 15 3
257 196
257 205
327 205
2 0 4 0 0 0 0 8 0 0 18 2
257 160
257 137
2 0 2 0 0 0 0 4 0 0 14 3
365 212
365 258
327 258
1 1 2 0 0 0 0 1 5 0 0 2
327 278
327 241
2 2 9 0 0 0 0 5 3 0 0 2
327 221
327 160
1 0 3 0 0 0 0 4 0 0 17 2
365 195
365 137
3 1 3 0 0 4224 0 3 6 0 0 2
345 137
465 137
1 1 4 0 0 4224 0 7 3 0 0 2
214 137
309 137
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 4
385 122 418 137
385 122 418 137
4 vout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 3
269 122 295 137
269 122 295 137
3 vin
-16 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 17
240 35 420 64
244 39 414 58
17 Voltage Regulator
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 23
546 48 682 92
550 52 678 84
23 Output
(+6V regulated)
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 25
11 49 171 93
15 53 167 85
25 Input
(+12V unregulated)
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 199
18 154 178 398
22 158 174 350
199 External Input 
Signal--A 200mV 
sine wave on a 
+12VDC signal 
produces our 
unregulated input 
voltage for 
simulation 
purposes only. 
This device is 
excluded from the 
PCB.
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 228
584 118 740 382
589 123 737 331
228 External 
Load--This is 
placed here for 
simulation 
purposes only. It 
is not part of 
the PCB. If you 
double-click on 
this device, you 
will notice that 
the "Exclude From 
PCB" checkbox is 
checked.
-13 0 0 0 400 0 0 0 0 1 2 1 49
7 Courier
0 0 0 8
201 70 274 87
205 74 269 83
8 PC Board
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.266667 0.000333333 0.000333333
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
