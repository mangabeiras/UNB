CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
13 70 515 411
7 5.000 V
7 5.000 V
3 GND
13 70 515 411
9437184 0
0
0
0
0
0
0
18
13 Logic Switch~
5 36 249 0 2 3
0 2 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 36 223 0 2 3
0 3 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 37 196 0 2 3
0 4 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 89 119 0 2 3
0 13 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 90 95 0 2 3
0 15 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 91 71 0 2 3
0 17 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 93 47 0 2 3
0 19 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 42 107 0 2 3
0 14 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 42 81 0 2 3
0 16 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 43 58 0 2 3
0 18 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 43 35 0 2 3
0 20 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 238 25 0 2 3
0 21 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8903 0 0
0
0
13 Logic Switch~
5 361 27 0 2 3
0 22 -99
0
0 0 20592 0
2 5V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3834 0 0
0
0
9 CA 7-Seg~
184 410 75 0 18 19
10 20 19 18 17 16 15 14 13 22
0 0 0 0 0 0 0 0 1
0
0 0 20592 0
5 REDCA
16 -41 51 -33
0
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
3363 0 0
0
0
9 CC 7-Seg~
183 289 75 0 9 19
10 20 19 18 17 16 15 14 13 21
0
0 0 20592 0
5 REDCC
16 -41 51 -33
0
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
7668 0 0
0
0
14 Ascii Display~
172 329 241 0 42 43
0 6 7 8 9 10 11 12 5 0
48 21608 26995 8297 29472 24864 29797 29556 8224 28518
8308 26725 8268 17220 8224 8224 8224 25705 29552 27745
31008 25701 30313 25445 11822 8224 8224 8224 8224 8224
8224 8224 8224
0
0 0 20592 0
4 1MEG
-15 -42 13 -34
0
0
0
102 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
%DE %5 0 %V
%DF %6 0 %V
%DG %7 0 %V
%DH %8 0 %V
0
0
0
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
82 0 0 0 1 0 0 0
4 DISP
4718 0 0
0
0
10 StopLight~
181 97 223 0 3 7
0 4 3 2
0
0 0 20592 0
4 1MEG
-15 -42 13 -34
0
0
0
37 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
0
0
0
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
3 SEM
3874 0 0
0
0
10 Ascii Key~
169 210 174 0 11 11
0 12 11 10 9 8 7 6 5 0
0 46
0
0 0 20528 0
0
0
0
0
0
0
0
0
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
3 KBD
6671 0 0
0
0
38
1 3 2 0 0 4224 0 1 17 0 0 4
48 249
70 249
70 237
81 237
2 1 3 0 0 4224 0 17 2 0 0 2
81 223
48 223
1 1 4 0 0 4224 0 3 17 0 0 4
49 196
70 196
70 209
81 209
8 8 5 0 0 4224 0 18 16 0 0 3
189 198
189 272
257 272
1 7 6 0 0 4224 0 16 18 0 0 3
263 210
195 210
195 198
6 2 7 0 0 8320 0 18 16 0 0 3
201 198
201 219
263 219
3 5 8 0 0 4224 0 16 18 0 0 3
263 228
207 228
207 198
4 4 9 0 0 8320 0 18 16 0 0 3
213 198
213 237
263 237
5 3 10 0 0 8320 0 16 18 0 0 3
263 246
219 246
219 198
2 6 11 0 0 4224 0 18 16 0 0 3
225 198
225 255
263 255
7 1 12 0 0 8320 0 16 18 0 0 3
263 264
231 264
231 198
8 8 13 0 0 4160 0 14 0 0 20 2
431 111
431 129
7 7 14 0 0 4160 0 14 0 0 20 2
425 111
425 129
6 6 15 0 0 4160 0 14 0 0 20 2
419 111
419 129
5 5 16 0 0 4160 0 14 0 0 20 2
413 111
413 129
4 4 17 0 0 4160 0 14 0 0 20 2
407 111
407 129
3 3 18 0 0 4160 0 14 0 0 20 2
401 111
401 129
2 2 19 0 0 4160 0 14 0 0 20 2
395 111
395 129
1 1 20 0 0 4160 0 14 0 0 20 2
389 111
389 129
1 1 1 0 0 12448 0 0 0 0 0 4
150 14
154 14
154 129
456 129
1 8 13 0 0 4288 0 4 0 0 20 2
101 119
154 119
1 7 14 0 0 4288 0 8 0 0 20 2
54 107
154 107
1 6 15 0 0 4288 0 5 0 0 20 2
102 95
154 95
1 5 16 0 0 4288 0 9 0 0 20 2
54 81
154 81
1 4 17 0 0 4288 0 6 0 0 20 2
103 71
154 71
1 3 18 0 0 4288 0 10 0 0 20 2
55 58
154 58
1 2 19 0 0 4288 0 7 0 0 20 2
105 47
154 47
1 1 20 0 0 4288 0 11 0 0 20 2
55 35
154 35
8 8 13 0 0 64 0 15 0 0 20 2
310 111
310 129
7 7 14 0 0 64 0 15 0 0 20 2
304 111
304 129
6 6 15 0 0 64 0 15 0 0 20 2
298 111
298 129
5 5 16 0 0 64 0 15 0 0 20 2
292 111
292 129
4 4 17 0 0 64 0 15 0 0 20 2
286 111
286 129
3 3 18 0 0 64 0 15 0 0 20 2
280 111
280 129
2 2 19 0 0 64 0 15 0 0 20 2
274 111
274 129
1 1 20 0 0 64 0 15 0 0 20 2
268 111
268 129
9 1 21 0 0 8320 0 15 12 0 0 3
289 33
289 25
250 25
9 1 22 0 0 8320 0 14 13 0 0 3
410 39
410 27
373 27
0
0
17 0 0
0
0
3 Vin
-1.5 -0.7 0.01
3 Vcc
10 14 1
100 0 1 100000
0 0.0005 2.5e-006 2.5e-006 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
0.002 0 0.09 -0.09 0.002 0.002
16 0
0 0.0005 10
0
0 0 100 100 0 0
98 66 294 126
0 0 0 0
294 66
98 66
294 66
294 126
0 0
1e+007 1 12.16 12.184 1e+007 1e+007
12403 0
0 3e+006 5e+006
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
2000 1 2.38857 0 1999 1999
16 0
0 500 1000
0
0 0 100 100 0 0
98 66 296 126
0 0 0 0
296 66
98 66
296 66
296 126
0 0
1e+006 1 -3.55271e-015 0 999999 999999
12403 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
