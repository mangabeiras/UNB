CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 80 30 100 9
0 66 640 259
8  5.000 V
8  5.000 V
3 GND
4.9505 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 259
9961490 2
0
0
0
0
0
0
6
5 SAVE-
218 228 131 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
5 SAVE1
-11 -36 24 -28
0
0
20 *Combine
*TRAN 0 15
0
0
0
1

0 0
0 0 0 0 1 0 0 0
4 SAVE
8953 0 0
0
0
5 SAVE-
218 314 131 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
5 SAVE2
-11 -36 24 -28
0
0
20 *Combine
*TRAN 0 15
0
0
0
1

0 0
0 0 0 0 1 0 0 0
4 SAVE
4441 0 0
0
0
11 Signal Gen~
195 175 151 0 24 64
0 3 2 1 86 9 10 0 0 0
0 0 0 0 0 0 0 1063828016 0 1097859072
0 1065353216 869711765 869711765 1066192077
20
0 0.909091 0 15 0 1 1e-007 1e-007 1.1 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
5 0/15V
-17 -28 18 -20
2 V1
-7 -38 7 -30
0
0
43 %D %1 %2 DC 0 PULSE(0 15 0 1 100n 100n 1.1)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
7 Ground~
168 301 187 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
5 Fuse~
219 273 131 0 2 5
0 3 4
5 Fuse~
0 0 4928 0
5 500mA
-17 -16 18 -8
2 F1
-7 -26 7 -18
0
0
11 %D %1 %2 %S
0
26 alias:XFUSE {CURRENT=500m}
4 FUSE
5

0 1 2 1 2 0
88 0 0 0 1 0 0 0
1 F
5394 0 0
0
0
9 Resistor~
219 354 131 0 4 5
0 4 2 0 -1
9 Resistor~
0 0 864 0
2 10
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
7734 0 0
0
0
4
1 1 3 0 0 4224 0 5 3 0 0 4
251 131
214 131
214 146
206 146
2 1 4 0 0 4224 0 5 6 0 0 2
295 131
336 131
1 0 2 0 0 4096 0 4 0 0 4 2
301 181
301 156
2 2 2 0 0 12416 0 6 3 0 0 4
372 131
388 131
388 156
206 156
0
0
16 0 0
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 1.01 0.0275 0.0275
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2672 8550976 100 100 0 0
98 66 608 126
0 259 640 452
608 66
98 66
608 71
608 125
0 0
5.26396e-315 0 5.22127e-315 4.97973e-315 5.26396e-315 5.26396e-315
12409 0
4 0.3 10
1
339 131
0 4 0 0 1	6 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
