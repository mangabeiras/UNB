CircuitMaker Text
5.6
Probes: 2
V2_1
Transient Analysis
0 178 137 65280
U2_3
Transient Analysis
1 336 137 65535
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
245 80 857 634
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
2 4 0.500000 0.500000
245 357 857 634
12058626 0
0
6 Title:
5 Name:
0
0
0
9
7 Ground~
168 198 171 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3964 0 0
2
36626.4 0
0
7 Ground~
168 365 181 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5105 0 0
2
36626.4 1
0
7 Ground~
168 381 96 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3782 0 0
2
36626.4 2
0
2 +V
167 251 109 0 1 3
0 4
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3573 0 0
2
36626.4 3
0
11 Signal Gen~
195 134 141 0 19 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V2
-8 -40 6 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7479 0 0
2
36626.4 4
0
7 gain:A~
219 287 145 0 4 9
0 3 4 6 2
0
0 0 54096 0
4 GAIN
-5 -31 23 -23
2 U2
2 -41 16 -33
0
0
29 %D %%vd(%1,%2) %%vd(%3,%4) %M
0
9 type:gain
0
9

0 0 0 0 0 0 0 0 0 0
65 0 0 0 1 0 0 0
1 U
8839 0 0
2
36626.4 5
0
5 gain~
219 286 72 0 2 5
0 3 5
0
0 0 50000 0
4 GAIN
-7 -31 21 -23
2 U1
0 -41 14 -33
0
0
11 %D %1 %2 %M
0
9 type:gain
0
5

0 0 0 0 0 0
65 0 0 0 1 0 0 0
1 U
6131 0 0
2
36626.4 6
0
9 Resistor~
219 361 136 0 4 5
0 6 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6110 0 0
2
36626.4 7
0
9 Resistor~
219 356 72 0 4 5
0 5 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
9311 0 0
2
36626.4 8
0
9
1 2 2 0 0 8192 0 1 5 0 0 3
198 165
198 146
165 146
1 0 2 0 0 0 0 2 0 0 4 2
365 175
365 154
1 2 2 0 0 0 0 3 9 0 0 3
381 90
381 72
374 72
4 2 2 0 0 4224 0 6 8 0 0 4
325 154
387 154
387 136
379 136
1 0 3 0 0 8192 0 7 0 0 6 3
262 72
199 72
199 136
1 1 3 0 0 4224 0 6 5 0 0 2
263 136
165 136
1 2 4 0 0 4224 0 4 6 0 0 3
251 118
251 154
263 154
1 2 5 0 0 4224 0 9 7 0 0 2
338 72
324 72
1 3 6 0 0 4224 0 8 6 0 0 2
343 136
325 136
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
4036 1210432 100 100 0 0
0 0 0 0
0 66 161 136
0 0
0 0
0 0
0 0
217 65
0 0 0 0 0 0
12401 0
4 1 3
1
225 72
0 3 0 0 1	0 5 0 0
3476 8550464 100 100 0 0
77 66 977 246
0 403 1024 740
977 66
77 66
977 66
977 246
0 0
4.94359e-315 0 5.27183e-315 1.58818e-314 4.94359e-315 4.94359e-315
12401 0
4 0.001 3
1
221 136
0 3 0 0 1	0 6 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
