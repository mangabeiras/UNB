CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 452
7 5.000 V
7 5.000 V
3 GND
0 66 640 452
9437184 0
0
0
0
0
0
0
15
13 Piezo Buzzer~
174 425 278 0 2 5
10 8 2
0
0 0 4208 0
4 .1uF
10 -16 38 -8
0
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
2 BZ
8953 0 0
0
0
13 Piezo Buzzer~
174 416 124 0 2 5
10 11 2
0
0 0 4208 0
4 .1uF
10 -16 38 -8
0
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
2 BZ
4441 0 0
0
0
12 SPST Switch~
165 424 236 0 2 5
0 3 8
0
0 0 20592 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3618 0 0
0
0
2 +V
167 460 217 0 1 3
0 3
0
0 0 53488 0
3 10V
12 -2 33 6
0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
11 SPDT Relay~
176 372 296 0 10 11
0 8 8 12 8 2 0 0 0 0
1
0
0 0 20592 0
7 12VSPDT
11 8 60 16
0
0
0
20 %D %1 %2 %3 %4 %5 %S
0
45 alias:XSPDTRELAY {PULLIN=9.6 RESISTANCE=1000}
4 DIP4
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 512 1 0 0 0
3 RLY
5394 0 0
0
0
7 Window~
179 284 241 0 4 9
0 8 13 8 14
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
7734 0 0
0
0
7 Window~
179 175 241 0 4 9
0 8 15 8 16
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
9914 0 0
0
0
7 Window~
179 62 239 0 4 9
0 8 17 8 18
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
3747 0 0
0
0
12 SPST Switch~
165 412 34 0 2 5
0 9 10
0
0 0 20592 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3549 0 0
0
0
7 Ground~
168 456 149 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
2 +V
167 454 16 0 1 3
0 9
0
0 0 53488 0
3 10V
12 -2 33 6
0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
7 Window~
179 280 79 0 4 9
0 11 10 19 20
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
8903 0 0
0
0
7 Window~
179 170 80 0 4 9
0 11 10 21 22
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
3834 0 0
0
0
7 Window~
179 59 81 0 4 9
0 11 10 23 24
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 WND
3363 0 0
0
0
7 Ground~
168 461 333 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
17
2 1 2 0 0 8192 0 1 15 0 0 3
456 278
461 278
461 327
2 1 2 0 0 0 0 2 10 0 0 3
447 124
456 124
456 143
5 0 2 0 0 8320 0 5 0 0 1 3
356 315
356 322
461 322
1 1 3 0 0 4224 0 3 4 0 0 3
441 236
460 236
460 226
3 4 8 0 0 12416 4 8 5 0 0 4
108 266
117 266
117 291
356 291
3 1 8 0 0 12416 5 7 8 0 0 6
221 268
230 268
230 282
128 282
128 257
108 257
3 1 8 0 0 12416 6 6 7 0 0 6
330 268
335 268
335 282
239 282
239 259
221 259
1 0 8 0 0 4224 7 6 0 0 9 2
330 259
391 259
2 2 8 0 0 0 7 5 3 0 0 4
386 271
391 271
391 236
407 236
1 1 8 0 0 4224 0 1 5 0 0 2
394 278
386 278
1 1 9 0 0 4224 0 9 11 0 0 3
429 34
454 34
454 25
2 2 10 0 0 4224 0 9 14 0 0 4
395 34
110 34
110 90
105 90
2 0 10 0 0 0 0 12 0 0 12 3
326 88
337 88
337 34
2 0 10 0 0 0 0 13 0 0 12 3
216 89
230 89
230 34
1 0 11 0 0 8192 0 13 0 0 17 3
216 98
238 98
238 124
1 0 11 0 0 8192 0 12 0 0 17 3
326 97
343 97
343 124
1 1 11 0 0 12416 0 14 2 0 0 4
105 99
120 99
120 124
385 124
4
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 44
29 128 350 155
33 132 340 151
44 Normally-Open Parallel Circuit Burgler Alarm
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 13
390 37 457 87
394 41 447 79
13 Enable
Alarm
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 13
398 181 465 231
402 185 455 223
13 Enable
Alarm
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 44
33 295 355 322
37 299 345 318
44 Normally-Closed Series Circuit Burgler Alarm
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 100 100 0 0
77 66 617 126
0 0 0 0
617 66
77 66
617 66
617 126
0 0
0.0005 0 1.2 -1.2 0.0005 0.0005
16 0
0 0.0001 10
0
0 0 100 100 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 -1.#IND -1.#IND 0 0
0 0
0 0.0002 10
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
