CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
0 66 640 259
144179216 0
0
0
0
0
0
0
8
5 SAVE-
218 130 22 0 64 64
0 0 0 0 0 0 0 0 0 0
1 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -1610612472
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
14 *DC 6.65 153 0
0
0
0
1

0 0
0 0 0 0 1 0 0 0
4 SAVE
8953 0 0
0
0
7 Ground~
168 62 163 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 239 141 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
9 V Source~
197 130 40 0 2 5
0 5 3
0
0 0 16736 0
2 0V
15 -2 29 6
2 V1
15 -12 29 -4
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
6153 0 0
0
0
9 V Source~
197 239 95 0 2 5
0 5 2
0
0 0 16992 0
3 10V
12 -2 33 6
3 VDS
12 -12 33 -4
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
5394 0 0
0
0
9 V Source~
197 62 127 0 2 5
0 4 2
0
0 0 16992 0
3 10V
12 -2 33 6
3 VGS
12 -12 33 -4
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
7734 0 0
0
0
7 Ground~
168 130 135 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
12 N-EMOS 3T:A~
219 124 93 0 3 7
0 3 4 2
12 N-EMOS 3T:A~
0 0 832 0
8 Si3454DV
18 0 74 8
2 Q1
39 -10 53 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TSOP-6
7

0 1 2 3 1 2 3 0
77 0 546 256 0 0 0 0
1 Q
3747 0 0
0
0
6
2 1 2 0 0 4224 0 5 3 0 0 2
239 116
239 135
1 2 3 0 0 4224 0 8 4 0 0 2
130 75
130 61
1 2 4 0 0 8320 0 6 8 0 0 3
62 106
62 102
106 102
1 2 2 0 0 0 0 2 6 0 0 2
62 157
62 148
1 1 5 0 0 8320 0 4 5 0 0 4
130 19
130 12
239 12
239 74
3 1 2 0 0 0 0 8 7 0 0 2
130 111
130 129
0
0
4 0 0
0
0
3 VDS
0.5 20 0.1
3 VGS
5 10 1
3 0 1 4
0 8e-007 1e-008 1e-008 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
3284 2259008 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
5.43943e-315 5.2221e-315 5.5705e-315 0 5.43813e-315 5.43813e-315
16 0
4 5 100
1
130 22
0 5 0 0 1	4 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
