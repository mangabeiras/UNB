CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 431
7 5.000 V
7 5.000 V
3 GND
0 66 640 431
9961472 0
0
0
0
0
0
0
12
5 SAVE-
218 215 121 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
12 *TRAN 0 5.04
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
7 Ground~
168 72 305 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
7 Ground~
168 215 296 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
10 Capacitor~
219 72 267 0 2 64
0 2 3
10 Capacitor~
0 0 848 90
4 22pF
8 5 36 13
2 C2
15 -5 29 3
0
0
18 %D %1 %2 %V IC=2.5
0
0
0
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
7 Ground~
168 147 161 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
2 +V
167 147 31 0 1 64
0 6
0
0 0 54128 0
2 5V
-5 -13 9 -5
3 VDD
-8 -23 13 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
12 N-MOSFET 3T~
219 137 131 0 3 64
0 5 3 2
12 N-MOSFET 3T~
0 0 848 0
4 NMOS
23 -4 51 4
2 M1
30 -14 44 -6
0
0
29 %D %1 %2 %3 %3 %M W=40U L=10U
0
0
0
7

0 1 2 3 1 2 3 -33686019
77 0 0 0 1 0 0 0
1 Q
9914 0 0
0
0
12 P-MOSFET 3T~
219 137 78 0 3 64
0 5 3 6
12 P-MOSFET 3T~
0 0 848 692
4 PMOS
23 -4 51 4
2 M2
30 -14 44 -6
0
0
29 %D %1 %2 %3 %3 %M W=80U L=10U
0
0
0
7

0 1 2 3 1 2 3 -33686019
109 0 0 0 1 0 0 0
1 Q
3747 0 0
0
0
8 Crystal~
219 147 241 0 2 64
0 3 4
8 Crystal~
0 0 848 0
9 3.5795MHZ
-29 -19 34 -11
4 XTAL
-12 -30 16 -22
0
0
11 %D %1 %2 %S
0
45 alias:XCRYSTAL {FREQ=3.58E6 RS=160 C=1.8E-11}
4 HC49
5

0 1 2 1 2 -33686019
88 0 0 0 0 0 0 0
4 XTAL
3549 0 0
0
0
10 Capacitor~
219 215 262 0 2 64
0 2 4
10 Capacitor~
0 0 848 90
4 22pF
9 4 37 12
2 C1
16 -6 30 2
0
0
18 %D %1 %2 %V IC=2.5
0
0
0
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
7931 0 0
0
0
9 Resistor~
219 215 170 0 2 64
0 4 5
9 Resistor~
0 0 4976 90
3 10k
5 6 26 14
2 RL
8 -4 22 4
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 150 202 0 2 64
0 3 4
9 Resistor~
0 0 880 0
4 220k
-14 -12 14 -4
2 RP
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
13
1 0 3 0 0 4096 0 12 0 0 8 2
132 202
72 202
2 0 4 0 0 4096 0 12 0 0 5 2
168 202
215 202
1 0 3 0 0 4096 0 9 0 0 8 2
136 241
72 241
2 0 4 0 0 4096 0 9 0 0 5 2
158 241
215 241
1 2 4 0 0 4224 0 11 10 0 0 2
215 188
215 253
1 1 2 0 0 4096 0 10 3 0 0 2
215 271
215 290
1 1 2 0 0 4224 0 4 2 0 0 4
72 276
72 302
72 302
72 299
0 2 3 0 0 8320 0 0 4 11 0 3
107 102
72 102
72 258
3 1 2 0 0 0 0 7 5 0 0 2
147 146
147 155
2 0 5 0 0 8320 0 11 0 0 12 3
215 152
215 100
147 100
2 2 3 0 0 0 0 8 7 0 0 4
127 63
107 63
107 140
127 140
1 1 5 0 0 0 0 8 7 0 0 2
147 90
147 113
3 1 6 0 0 4224 0 8 6 0 0 2
147 57
147 40
0
0
16 2 0
0
0
0
0 0 0
0
0 0 0
0 0 1 2
1e-005 1.1e-005 2e-008 2e-008 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
2296 8550464 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
1.1e-005 1.00056e-005 1.1e-005 1.00056e-005 9.944e-007 9.944e-007
0 0
4 3e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
