CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
6000.24 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 259
9961474 0
0
0
0
0
0
0
16
10 Capacitor~
219 122 75 0 2 64
0 8 5
10 Capacitor~
0 0 320 0
5 .01uF
-18 -18 17 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
8953 0 0
0
0
7 Ground~
168 313 118 0 1 64
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 69 108 0 1 64
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
2 +V
167 120 8 0 1 64
0 3
0
0 0 53600 90
4 +15V
-33 -6 -5 2
2 V1
-7 -15 7 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
5 SAVE-
218 298 52 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
26 *Combine
*TRAN -502m 492m
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SAVE-
218 76 75 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
26 *Combine
*TRAN -502m 492m
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
11 Signal Gen~
195 27 80 0 19 64
0 8 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1169915904 0 1047904911
20
1 6000 0 0.24 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 64 0
11 -240m/240mV
-39 -20 38 -12
2 V2
-7 -30 7 -22
0
0
39 %D %1 %2 DC 0 SIN(0 240m 6k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
7 Ground~
168 216 155 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
10 NPN Trans~
219 209 75 0 3 64
0 4 5 6
10 NPN Trans~
0 0 320 0
7 2N2222A
8 0 57 8
2 Q1
25 -10 39 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 -33686019
81 0 0 0 1 0 0 0
1 Q
3549 0 0
0
0
10 Capacitor~
219 259 126 0 2 64
0 2 6
10 Capacitor~
0 0 320 90
5 .01uF
11 0 46 8
2 C2
22 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
7931 0 0
0
0
10 Capacitor~
219 265 52 0 2 64
0 4 7
10 Capacitor~
0 0 320 0
5 .01uF
-18 -18 17 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
9325 0 0
0
0
9 Resistor~
219 216 28 0 3 64
0 3 4 1
9 Resistor~
0 0 4448 270
3 675
7 0 28 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 147 27 0 3 64
0 3 5 1
9 Resistor~
0 0 4448 270
3 18k
7 0 28 8
2 R2
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.3
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 313 80 0 3 64
0 2 7 -1
9 Resistor~
0 0 4448 90
3 10K
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 216 123 0 3 64
0 2 6 -1
9 Resistor~
0 0 352 90
3 200
7 0 28 8
2 R4
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 147 122 0 3 64
0 2 5 -1
9 Resistor~
0 0 352 90
4 3.3k
8 0 36 8
2 R5
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
4718 0 0
0
0
16
1 0 3 0 0 4096 0 4 0 0 9 2
131 6
147 6
1 0 4 0 0 4224 0 11 0 0 14 2
256 52
216 52
2 2 5 0 0 4224 0 1 9 0 0 2
131 75
203 75
1 1 2 0 0 4096 0 14 2 0 0 2
313 98
313 112
2 1 2 0 0 8192 0 7 3 0 0 3
58 85
69 85
69 102
0 1 2 0 0 0 0 0 15 8 0 2
216 147
216 141
1 0 2 0 0 0 0 8 0 0 8 4
216 149
216 151
216 151
216 147
1 1 2 0 0 8320 0 16 10 0 0 4
147 140
147 147
259 147
259 135
1 1 3 0 0 8320 0 13 12 0 0 4
147 9
147 6
216 6
216 10
0 2 5 0 0 0 0 0 13 3 0 2
147 75
147 45
2 0 6 0 0 8320 0 10 0 0 13 3
259 117
259 98
216 98
2 0 5 0 0 0 0 16 0 0 3 2
147 104
147 75
3 2 6 0 0 0 0 9 15 0 0 2
216 93
216 105
1 2 4 0 0 0 0 9 12 0 0 2
216 57
216 46
2 2 7 0 0 4224 0 11 14 0 0 3
274 52
313 52
313 62
1 1 8 0 0 4224 0 1 7 0 0 2
113 75
58 75
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
100 0 1 1e+006
0 0.0008333 4.167e-006 4.167e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3852 8550464 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
4.83693e-315 0 5.23039e-315 1.58404e-314 4.83693e-315 4.83693e-315
16 0
4 0.0002 10
2
84 75
0 8 0 0 1	0 16 0 0
300 52
0 7 0 0 1	0 15 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
