CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 3
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
0 66 640 259
12058626 0
0
0
0
0
0
0
12
5 SAVE-
218 306 42 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 D
3 -26 10 -18
0
0
0
16 *TRAN -4.43 4.43
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 91 42 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 C
3 -26 10 -18
0
0
0
26 *Combine
*TRAN -5.43 5.43
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SAVE-
218 206 69 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
26 *Combine
*TRAN -5.43 5.43
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SAVE-
218 211 42 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
26 *Combine
*TRAN -5.43 5.43
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
7 Ground~
168 312 124 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 78 139 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7734 0 0
0
0
11 Signal Gen~
195 38 47 0 19 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 16704 0
5 -1/1V
-17 -28 18 -20
2 V1
-7 -38 7 -30
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
8 V-Math1~
219 166 42 0 2 5
0 6 5
8 V-Math1~
0 0 5184 0
6 UNARYV
-21 -26 21 -18
2 M1
-7 -36 7 -28
4 -(V)
-13 -14 15 -6
0
11 %D %1 %2 %S
0
0
4 -(V)
5

0 1 2 1 2 0
88 0 0 0 0 0 0 0
1 M
3747 0 0
0
0
8 V-Math1~
219 165 74 0 2 5
0 6 4
8 V-Math1~
0 0 5184 0
6 ATANHV
-21 -26 21 -18
2 M2
-7 -36 7 -28
8 ATANH(V)
-27 -14 29 -6
0
11 %D %1 %2 %S
0
0
8 ATANH(V)
5

0 1 2 1 2 0
88 0 0 0 0 0 0 0
1 M
3549 0 0
0
0
8 V-Math2~
219 264 51 0 3 7
0 5 4 3
8 V-Math2~
0 0 5184 0
4 ADDV
-14 -36 14 -27
2 M3
-7 -46 7 -38
6 V(A+B)
-20 -23 22 -15
0
14 %D %1 %2 %3 %S
0
0
6 V(A+B)
7

0 1 2 3 1 2 3 0
88 0 0 256 0 0 0 0
1 M
7931 0 0
0
0
9 Resistor~
219 312 85 0 3 5
0 2 3 -1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 105 99 0 3 5
0 2 6 -1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
8903 0 0
0
0
9
1 1 2 0 0 4096 0 11 5 0 0 2
312 103
312 118
3 2 3 0 0 8320 0 10 11 0 0 3
298 42
312 42
312 67
2 2 4 0 0 12416 0 9 10 0 0 4
199 74
205 74
205 51
230 51
2 1 5 0 0 4224 0 8 10 0 0 2
200 42
230 42
1 0 6 0 0 4096 0 9 0 0 6 2
131 74
105 74
2 0 6 0 0 4096 0 12 0 0 7 2
105 81
105 42
1 1 6 0 0 4224 0 7 8 0 0 2
69 42
132 42
1 0 2 0 0 8192 0 12 0 0 9 3
105 117
105 122
78 122
2 1 2 0 0 8320 0 7 6 0 0 3
69 52
78 52
78 133
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 0.005 5e-006 5e-006 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
860 8550464 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
4.94359e-315 0 5.36716e-315 1.59771e-314 4.94359e-315 5.4086e-315
16 0
4 0.001 3
1
312 51
0 3 0 0 2	0 2 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
