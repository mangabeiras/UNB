CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 300 100 9
0 66 572 394
7 5.000 V
7 5.000 V
3 GND
3125 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 572 394
9961474 0
0
0
0
0
0
0
21
5 SAVE-
218 275 91 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
20 *Combine
*TRAN 0 10
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
9 Terminal~
194 334 92 0 1 64
0 3
0
0 0 53568 26894
6 Output
-24 -18 18 -10
2 T1
-10 -26 4 -18
0
0
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
1 T
4441 0 0
0
0
7 Ground~
168 247 197 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
2 +V
167 128 199 0 1 64
0 4
0
0 0 53600 -19276
3 -5V
-12 2 9 10
2 V1
-9 -8 5 0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
7 Ground~
168 128 270 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
11 Signal Gen~
195 81 244 0 24 64
0 8 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1148846080 1092616192 0
953267991 869711765 869711765 973279855 981668463
20
0 1000 10 0 0.0001 1e-007 1e-007 0.0005 0.001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 320 0
5 10/0V
-17 -28 18 -20
2 V2
-7 -38 7 -30
0
0
48 %D %1 %2 DC 0 PULSE(10 0 100u 100n 100n 500u 1m)
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
7 Ground~
168 81 168 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
2 +V
167 166 16 0 1 64
0 9
0
0 0 53600 0
4 +10V
-13 -13 15 -5
2 V3
-7 -26 7 -18
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
12 NPN Trans:C~
219 242 130 0 3 64
0 3 6 7
12 NPN Trans:C~
0 0 320 0
6 2N3904
10 13 52 21
2 Q1
34 -14 48 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 0 0 0
1 Q
3549 0 0
0
0
12 NPN Trans:C~
219 90 130 0 3 64
0 10 11 2
12 NPN Trans:C~
0 0 320 512
6 2N3904
-56 13 -14 21
2 Q2
-56 -15 -42 -7
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 0 0 0
1 Q
7931 0 0
0
0
10 Capacitor~
219 114 104 0 2 64
0 10 6
10 Capacitor~
0 0 320 0
5 .02uF
-18 -18 17 -10
2 C1
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
9325 0 0
0
0
10 Capacitor~
219 216 80 0 2 64
0 11 3
10 Capacitor~
0 0 320 0
5 100pF
-17 -19 18 -11
2 C2
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
8903 0 0
0
0
6 Diode~
219 198 172 0 2 64
0 6 5
6 Diode~
0 0 320 26894
5 1N914
-48 -3 -13 5
2 D1
23 -12 37 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
3834 0 0
0
0
6 Diode~
219 247 172 0 2 64
0 7 2
6 Diode~
0 0 320 26894
5 1N914
14 -4 49 4
2 D2
24 -12 38 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
3363 0 0
0
0
10 Capacitor~
219 153 239 0 2 64
0 8 5
10 Capacitor~
0 0 320 0
5 100pF
-14 -19 21 -11
2 C3
-4 -29 10 -21
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
7668 0 0
0
0
9 Resistor~
219 81 54 0 4 64
0 10 9 0 1
9 Resistor~
0 0 352 90
2 1k
-22 -4 -8 4
2 R1
7 -12 21 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 247 55 0 4 64
0 3 9 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R2
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 217 103 0 2 64
0 3 11
9 Resistor~
0 0 352 180
3 47k
-11 -11 10 -3
2 R3
10 -12 24 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 128 154 0 3 64
0 4 11 1
9 Resistor~
0 0 352 90
4 470k
5 -3 33 5
2 R4
12 -13 26 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 310 125 0 2 64
0 5 3
9 Resistor~
0 0 352 90
3 10k
-25 -4 -4 4
2 R5
-22 -14 -8 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 144 56 0 4 64
0 6 9 0 1
9 Resistor~
0 0 352 90
3 15k
6 -4 27 4
2 R6
9 -14 23 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
24
1 0 3 0 0 4096 0 2 0 0 14 2
322 91
310 91
1 1 4 0 0 4224 0 19 4 0 0 2
128 172
128 184
2 0 5 0 0 4096 0 13 0 0 8 2
198 182
198 239
1 0 6 0 0 4096 0 13 0 0 11 2
198 162
198 130
2 1 2 0 0 4096 0 14 3 0 0 2
247 182
247 191
3 1 7 0 0 4224 0 9 14 0 0 2
247 148
247 162
1 1 8 0 0 4224 0 15 6 0 0 2
144 239
112 239
1 2 5 0 0 8320 0 20 15 0 0 3
310 143
310 239
162 239
2 0 9 0 0 4096 0 21 0 0 24 2
144 38
144 32
1 0 6 0 0 0 0 21 0 0 11 2
144 74
144 104
2 2 6 0 0 12416 0 11 9 0 0 4
123 104
166 104
166 130
224 130
1 0 10 0 0 4096 0 11 0 0 22 2
105 104
81 104
2 1 2 0 0 4224 0 6 5 0 0 3
112 249
128 249
128 264
2 0 3 0 0 8320 0 20 0 0 21 3
310 107
310 91
247 91
2 0 11 0 0 4096 0 19 0 0 19 2
128 136
128 130
2 0 3 0 0 0 0 12 0 0 21 2
225 80
247 80
1 0 3 0 0 0 0 18 0 0 21 2
235 103
247 103
1 0 11 0 0 8192 0 12 0 0 19 3
207 80
188 80
188 103
2 2 11 0 0 4224 0 10 18 0 0 6
104 130
154 130
154 119
178 119
178 103
199 103
3 1 2 0 0 0 0 10 7 0 0 2
81 148
81 162
1 1 3 0 0 0 0 17 9 0 0 2
247 73
247 112
1 1 10 0 0 4224 0 16 10 0 0 2
81 72
81 112
1 0 9 0 0 4096 0 8 0 0 24 2
166 25
166 32
2 2 9 0 0 8320 0 16 17 0 0 4
81 36
81 32
247 32
247 37
2
-16 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 25
374 61 524 114
378 65 518 103
25 Monostable
Multivibrator
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 60
337 114 537 178
341 118 533 166
60 Triggers on the falling 
edge of the Signal Gen 
output.
0
16 0 1
0
0
0
0 0 0
0
0 0 0
200 0 1 1e+006
0 0.0016 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
