CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 300 100 9
0 66 640 452
7 5.000 V
7 5.000 V
3 GND
10000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 452
9961474 0
0
0
0
0
0
0
26
5 SAVE-
218 52 92 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
14 *TRAN 41m 10.5
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 264 91 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
14 *TRAN 41m 10.5
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
9 .NODESET~
208 291 71 0 1 64
0 3
0
0 0 53568 0
3 10V
-10 -15 11 -7
4 CMD1
-13 -25 15 -17
0
0
17 .NODESET V(%1)=%V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
3 CMD
3618 0 0
0
0
9 .NODESET~
208 37 72 0 1 64
0 4
0
0 0 53568 0
2 0V
-7 -15 7 -7
4 CMD2
-14 -25 14 -17
0
0
17 .NODESET V(%1)=%V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
3 CMD
6153 0 0
0
0
7 Ground~
168 166 283 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
11 Signal Gen~
195 107 264 0 24 64
0 6 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1176256512 0 1092616192
0 869711765 869711765 944879383 953267991
20
0 10000 0 10 0 1e-007 1e-007 5e-005 0.0001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 320 0
5 0/10V
-17 -28 18 -20
2 V1
-7 -38 7 -30
0
0
46 %D %1 %2 DC 0 PULSE(0 10 0 100n 100n 50u 100u)
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
2 +V
167 164 199 0 1 64
0 5
0
0 0 53600 180
4 -10V
-14 -1 14 7
2 V2
-7 -11 7 -3
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
7 Ground~
168 247 167 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
7 Ground~
168 81 168 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
2 +V
167 166 16 0 1 64
0 11
0
0 0 53600 0
4 +10V
-13 -13 15 -5
2 V3
-7 -26 7 -18
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
12 NPN Trans:C~
219 242 130 0 3 64
0 3 10 2
12 NPN Trans:C~
0 0 320 0
6 2N3904
10 13 52 21
2 Q1
34 -14 48 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 0 0 0
1 Q
9325 0 0
0
0
12 NPN Trans:C~
219 90 130 0 3 64
0 4 9 2
12 NPN Trans:C~
0 0 320 512
6 2N3904
-56 13 -14 21
2 Q2
-56 -15 -42 -7
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 0 0 0
1 Q
8903 0 0
0
0
10 Capacitor~
219 112 80 0 2 64
0 4 10
10 Capacitor~
0 0 320 0
5 200pF
-12 -20 23 -12
2 C1
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3834 0 0
0
0
10 Capacitor~
219 216 80 0 2 64
0 9 3
10 Capacitor~
0 0 320 0
5 200pF
-17 -19 18 -11
2 C2
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3363 0 0
0
0
6 Diode~
219 113 197 0 2 64
0 9 8
6 Diode~
0 0 320 26894
5 1N914
-48 -3 -13 5
2 D1
23 -12 37 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
7668 0 0
0
0
6 Diode~
219 215 197 0 2 64
0 10 7
6 Diode~
0 0 320 26894
5 1N914
14 -4 49 4
2 D2
24 -12 38 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
4718 0 0
0
0
10 Capacitor~
219 142 228 0 2 64
0 8 6
10 Capacitor~
0 0 320 0
5 200pF
-14 -17 21 -9
2 C3
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3874 0 0
0
0
10 Capacitor~
219 191 228 0 2 64
0 6 7
10 Capacitor~
0 0 320 0
5 200pF
-14 -17 21 -9
2 C4
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
6671 0 0
0
0
9 Resistor~
219 81 54 0 4 64
0 4 11 0 1
9 Resistor~
0 0 352 90
2 1k
-22 -4 -8 4
2 R1
7 -12 21 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 113 103 0 2 64
0 10 4
9 Resistor~
0 0 352 180
3 39k
-11 -12 10 -4
2 R2
9 -15 23 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 247 55 0 4 64
0 3 11 0 1
9 Resistor~
0 0 352 90
2 1k
8 -5 22 3
2 R3
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 217 103 0 2 64
0 3 9
9 Resistor~
0 0 352 180
3 39k
-11 -11 10 -3
2 R4
10 -12 24 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 128 154 0 3 64
0 5 9 1
9 Resistor~
0 0 352 90
4 390k
5 -3 33 5
2 R5
12 -13 26 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 200 154 0 3 64
0 5 10 1
9 Resistor~
0 0 352 90
4 390k
-32 -3 -4 5
2 R6
-25 -13 -11 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 303 116 0 2 64
0 7 3
9 Resistor~
0 0 352 90
3 10k
-25 -4 -4 4
2 R7
-22 -14 -8 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
9 Resistor~
219 22 122 0 2 64
0 8 4
9 Resistor~
0 0 352 90
3 10k
6 -5 27 3
2 R8
9 -15 23 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
31
1 0 3 0 0 4096 0 3 0 0 11 2
291 83
291 91
1 0 4 0 0 4096 0 4 0 0 12 2
37 84
37 92
1 0 5 0 0 4096 0 7 0 0 15 2
164 184
164 178
2 1 2 0 0 4224 0 6 5 0 0 3
138 269
166 269
166 277
1 0 6 0 0 8320 0 6 0 0 8 3
138 259
166 259
166 228
2 0 7 0 0 4096 0 16 0 0 9 2
215 207
215 228
2 0 8 0 0 4096 0 15 0 0 10 2
113 207
113 228
2 1 6 0 0 0 0 17 18 0 0 2
151 228
182 228
1 2 7 0 0 8320 0 25 18 0 0 3
303 134
303 228
200 228
1 1 8 0 0 8320 0 26 17 0 0 3
22 140
22 228
133 228
2 0 3 0 0 8320 0 25 0 0 28 3
303 98
303 91
247 91
2 0 4 0 0 8320 0 26 0 0 29 3
22 104
22 92
81 92
1 0 9 0 0 4224 0 15 0 0 24 2
113 187
113 130
1 0 10 0 0 4224 0 16 0 0 25 2
215 187
215 130
1 1 5 0 0 8320 0 23 24 0 0 4
128 172
128 178
200 178
200 172
2 0 9 0 0 0 0 23 0 0 24 2
128 136
128 130
2 0 10 0 0 0 0 24 0 0 25 2
200 136
200 130
2 0 3 0 0 0 0 14 0 0 28 2
225 80
247 80
1 0 3 0 0 0 0 22 0 0 28 2
235 103
247 103
1 0 9 0 0 0 0 14 0 0 24 3
207 80
188 80
188 103
2 0 10 0 0 0 0 13 0 0 25 3
121 80
145 80
145 103
1 0 4 0 0 0 0 13 0 0 29 2
103 80
81 80
2 0 4 0 0 0 0 20 0 0 29 2
95 103
81 103
2 2 9 0 0 0 0 12 22 0 0 6
104 130
154 130
154 120
181 120
181 103
199 103
2 1 10 0 0 0 0 11 20 0 0 6
224 130
173 130
173 113
154 113
154 103
131 103
3 1 2 0 0 0 0 12 9 0 0 2
81 148
81 162
3 1 2 0 0 0 0 11 8 0 0 2
247 148
247 161
1 1 3 0 0 0 0 21 11 0 0 2
247 73
247 112
1 1 4 0 0 0 0 19 12 0 0 2
81 72
81 112
1 0 11 0 0 4096 0 10 0 0 31 2
166 25
166 32
2 2 11 0 0 8320 0 19 21 0 0 4
81 36
81 32
247 32
247 37
2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 155
340 77 540 221
344 81 536 193
155 Since this is a 
symetrical bistable 
circuit, the nodeset 
(.NS) devices are used 
to help the simulation 
converge into two 
distinct states.
-16 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 23
341 18 491 71
345 22 485 60
23 Bistable
Multivibrator
0
16 0 1
0
0
0
0 0 0
0
0 0 0
200 0 1 1e+006
0 0.0005 2e-006 2e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
896 8550464 100 100 0 0
77 66 977 276
0 401 1024 742
977 66
77 66
977 66
977 276
0 0
4.94359e-315 0 5.30706e-315 1.5917e-314 4.94359e-315 4.94359e-315
16 0
4 0.0001 10
1
215 163
0 10 0 0 1	0 14 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
