CircuitMaker Text
5.6
Probes: 5
CMD1_1
AC Analysis
0 288 122 65280
CMD1_1
DC Sweep
0 288 122 65280
CMD1_1
Operating Point
0 288 122 65280
CMD1_1
Fourier Analysis
0 288 122 65280
out
Transient Analysis
0 276 120 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
231 152 911 669
7 5.000 V
7 5.000 V
3 GND
2000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
2 4 0.500000 0.500000
231 411 911 669
12058624 0
0
0
0
0
0
0
17
4 .IC~
207 237 68 0 1 64
0 3
0
0 0 53584 0
2 2V
-7 -16 7 -8
4 CMD1
-14 -26 14 -18
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
3 CMD
3760 0 0
2
36626.6 0
0
4 .IC~
207 74 105 0 1 64
0 5
0
0 0 53584 0
2 0V
-7 -16 7 -8
4 CMD2
-14 -26 14 -18
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
3 CMD
5673 0 0
2
36626.6 1
0
7 Ground~
168 126 256 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3256 0 0
2
36626.6 3
0
7 Ground~
168 66 197 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3672 0 0
2
36626.6 4
0
7 Ground~
168 27 201 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
6260 0 0
2
36626.6 5
0
2 +V
167 151 166 0 1 64
0 7
0
0 0 54128 -19276
4 -12V
-13 10 15 18
2 V1
-6 0 8 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
7667 0 0
2
36626.6 6
0
2 +V
167 151 87 0 1 64
0 8
0
0 0 54128 0
4 +12V
-14 -14 14 -6
2 V2
-7 -24 7 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3778 0 0
2
36626.6 7
0
10 Capacitor~
219 186 44 0 2 64
0 9 3
10 Capacitor~
0 0 848 0
6 0.01uF
-21 -18 21 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
9961 0 0
2
36626.6 8
0
8 Op-Amp5~
219 151 122 0 5 64
0 5 4 8 7 3
8 Op-Amp5~
0 0 848 0
5 UA741
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 -33686019
88 -1 258 0 1 0 0 0
1 U
6573 0 0
2
36626.6 9
0
10 Capacitor~
219 66 166 0 2 64
0 2 5
10 Capacitor~
0 0 848 90
6 0.01uf
12 0 54 8
2 C2
26 -10 40 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
8204 0 0
2
36626.6 10
0
13 Var Resistor~
219 262 210 0 3 64
0 4 4 6
13 Var Resistor~
0 0 848 90
7 50k 60%
12 -3 61 5
2 R1
26 -15 40 -7
0
0
32 %DA %1 %2 30000
%DB %2 %3 20000
0
0
4 SIP3
7

0 1 2 3 1 2 3 -33686019
82 0 272 0 1 0 0 0
1 R
961 0 0
2
36626.6 11
0
6 Diode~
219 211 151 0 2 64
0 6 3
6 Diode~
0 0 848 90
5 1N914
11 0 46 8
2 D1
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.7
5

0 1 2 1 2 -33686019
68 -1 280 0 1 0 0 0
1 D
4687 0 0
2
36626.6 12
0
6 Diode~
219 313 148 0 2 64
0 3 6
6 Diode~
0 0 848 26894
5 1N914
11 0 46 8
2 D2
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.7
5

0 1 2 1 2 -33686019
68 -1 280 0 1 0 0 0
1 D
7852 0 0
2
36626.6 13
0
9 Resistor~
219 117 44 0 2 64
0 5 9
9 Resistor~
0 0 880 0
3 12K
-11 -14 10 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3222 0 0
2
36626.6 14
0
9 Resistor~
219 27 167 0 3 64
0 2 5 -1
9 Resistor~
0 0 880 90
3 12k
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
496 0 0
2
36626.6 15
0
9 Resistor~
219 126 219 0 3 64
0 2 4 -1
9 Resistor~
0 0 880 90
3 12k
7 0 28 8
2 R4
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
8742 0 0
2
36626.6 16
0
9 Resistor~
219 266 151 0 2 64
0 6 3
9 Resistor~
0 0 880 90
3 12k
7 0 28 8
2 R5
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
4405 0 0
2
36626.6 17
0
21
1 0 3 0 0 8192 0 1 0 0 8 3
237 80
237 87
211 87
2 0 4 0 0 4096 0 11 0 0 3 2
254 208
236 208
1 0 4 0 0 16512 0 11 0 0 15 5
266 224
266 236
236 236
236 188
126 188
1 0 5 0 0 4096 0 2 0 0 14 2
74 117
74 128
2 0 6 0 0 8192 0 13 0 0 16 3
313 158
313 174
266 174
1 0 6 0 0 8320 0 12 0 0 16 3
211 161
211 174
266 174
2 0 3 0 0 0 0 12 0 0 10 2
211 141
211 122
2 0 3 0 0 8192 0 8 0 0 10 3
195 44
211 44
211 122
2 0 3 0 0 0 0 17 0 0 10 2
266 133
266 122
5 1 3 0 0 4224 0 9 13 0 0 3
169 122
313 122
313 138
4 1 7 0 0 4224 0 9 6 0 0 2
151 135
151 151
1 3 8 0 0 4224 0 7 9 0 0 2
151 96
151 109
2 0 5 0 0 4096 0 10 0 0 14 2
66 157
66 128
1 0 5 0 0 4224 0 9 0 0 20 2
133 128
27 128
2 2 4 0 0 0 0 9 16 0 0 3
133 116
126 116
126 201
1 3 6 0 0 0 0 17 11 0 0 2
266 169
266 188
1 1 2 0 0 4096 0 16 3 0 0 2
126 237
126 250
1 1 2 0 0 4224 0 10 4 0 0 2
66 175
66 191
1 1 2 0 0 0 0 15 5 0 0 2
27 185
27 195
1 2 5 0 0 0 0 14 15 0 0 3
99 44
27 44
27 149
1 2 9 0 0 4224 0 8 14 0 0 2
177 44
135 44
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 3
231 106 258 122
231 106 258 122
3 out
-16 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 22
357 9 587 38
361 13 581 32
22 Wien-Bridge Oscillator
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 442
356 31 628 315
360 35 624 259
442 The series and parallel RC 
networks (R2+C1 and R3+C2)in 
this circuit determine its 
oscillating frequency. The 
value of R1 sets the circuits 
gain. If the gain is close to 3 
(R1=2*R4) a sine wave will be 
produced. If the gain is 
greater than 3, the output will 
begin to clip. If the gain is 
less than 3, oscillation die 
out. Try using the script STEP 
VALUE function to vary R1 and 
view the output results.
33 .OPTIONS METHOD=GEAR ITL4=40.00

16 0 1
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 0.0025 1e-05 1e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
