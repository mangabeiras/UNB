CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 65 640 452
7 5.000 V
7 5.000 V
3 GND
0 65 640 452
9437184 0
0
0
0
0
0
0
19
7 74LS139
118 300 65 0 14 29
0 22 8 2 23 9 2 33 32 15
30 16 24 17 20
0
0 0 12528 0
7 74LS139
-24 -51 25 -43
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
13 type: digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 -33686019
65 0 0 0 1 1 0 0
1 U
8953 0 0
0
0
6 74LS75
103 173 74 0 14 29
0 28 27 21 26 25 21 22 34 8
35 23 36 9 37
0
0 0 12528 0
6 74LS75
-21 -51 21 -43
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
113 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 6 4 3 2 13 9 8 10
11 15 14 16 1 7 6 4 3 2
13 9 8 10 11 15 14 16 1 -33686019
65 0 0 512 1 1 0 0
1 U
4441 0 0
0
0
6 74LS93
109 80 56 0 8 17
0 2 2 21 25 28 27 26 25
0
0 0 12528 0
6 74LS93
-21 -35 21 -27
2 U5
-7 -45 7 -37
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 -33686019
65 0 0 0 1 1 0 0
1 U
3618 0 0
0
0
8 4-In OR~
219 566 159 0 5 21
0 18 12 11 10 3
0
0 0 112 0
4 4072
-14 -24 14 -16
3 U2A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 -33686019
65 0 0 0 2 1 3 0
1 U
6153 0 0
0
0
12 Hex Display~
7 327 153 0 4 9
10 7 6 5 4
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -52 17 -44
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5394 0 0
0
0
7 Ground~
168 249 125 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
12 2-In NOR:DM~
219 504 193 0 3 21
0 14 24 11
12 2-In NOR:DM~
0 0 112 0
6 74LS02
-21 -24 21 -16
3 U1D
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 4 2 0
1 U
9914 0 0
0
0
12 2-In NOR:DM~
219 504 230 0 3 21
0 13 16 10
12 2-In NOR:DM~
0 0 112 0
6 74LS02
-21 -24 21 -16
3 U1C
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 3 2 0
1 U
3747 0 0
0
0
12 2-In NOR:DM~
219 503 155 0 3 21
0 15 17 12
12 2-In NOR:DM~
0 0 112 0
6 74LS02
-21 -24 21 -16
3 U1B
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 2 2 0
1 U
3549 0 0
0
0
12 Quad D Flop~
47 278 219 0 9 19
0 9 23 8 22 7 6 5 4 3
0
0 0 4208 0
4 QDFF
-14 -44 14 -36
2 U6
-7 -54 7 -46
0
15 DVCC=16;DGND=8;
81 %D [%16bi %8bi %1i %2i %3i %4i %9i][%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 -33686019
65 0 0 0 1 1 0 0
1 U
7931 0 0
0
0
2 +V
167 484 287 0 1 3
0 29
0
0 0 53488 0
3 10V
12 -2 33 6
2 V1
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
7 Pulser~
4 40 137 0 9 9
0 38 39 21 40 0 0 5 5 2
0
0 0 20528 0
0
2 V2
-7 -38 7 -30
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8903 0 0
0
0
7 Ground~
168 13 78 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
11 4x4 Switch~
193 435 43 0 11 17
0 33 32 15 30 13 19 15 14 0
10 25
0
0 0 20592 0
0
3 SW1
-20 -52 1 -44
0
0
0
0
0
0
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
2 SW
3363 0 0
0
0
12 2-In NOR:DM~
219 502 117 0 3 21
0 19 20 18
12 2-In NOR:DM~
0 0 112 0
6 74LS02
-21 -24 21 -16
3 U1A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 2 0
1 U
7668 0 0
0
0
9 Resistor~
219 457 288 0 3 5
0 29 13 1
9 Resistor~
0 0 4208 90
2 1k
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 442 287 0 3 5
0 29 14 1
9 Resistor~
0 0 4208 90
2 1k
-7 -12 7 -4
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 428 287 0 3 5
0 29 15 1
9 Resistor~
0 0 4208 90
2 1k
-7 -12 7 -4
2 R3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 413 288 0 3 5
0 29 19 1
9 Resistor~
0 0 4208 90
2 1k
-7 -12 7 -4
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3789 0 0
0
0
49
5 9 3 0 0 12416 0 4 10 0 0 5
599 159
607 159
607 335
278 335
278 255
4 8 4 0 0 4224 0 5 10 0 0 3
318 177
318 225
302 225
3 7 5 0 0 4224 0 5 10 0 0 3
324 177
324 213
302 213
2 6 6 0 0 8320 0 5 10 0 0 3
330 177
330 201
302 201
1 5 7 0 0 8320 0 5 10 0 0 3
336 177
336 189
302 189
6 0 2 0 0 4096 0 1 0 0 7 2
262 101
249 101
3 1 2 0 0 8320 0 1 6 0 0 3
262 65
249 65
249 119
3 0 8 0 0 8320 0 10 0 0 27 3
254 213
223 213
223 65
1 0 9 0 0 8320 0 10 0 0 24 3
254 189
235 189
235 101
2 0 2 0 0 0 0 3 0 0 11 2
48 56
13 56
1 1 2 0 0 0 0 3 13 0 0 3
48 47
13 47
13 72
3 4 10 0 0 8320 0 8 4 0 0 4
525 230
544 230
544 173
549 173
3 3 11 0 0 8320 0 4 7 0 0 4
549 164
533 164
533 193
525 193
2 3 12 0 0 4224 0 4 9 0 0 2
549 155
524 155
1 0 13 0 0 4096 0 8 0 0 40 2
474 221
457 221
1 0 14 0 0 4096 0 7 0 0 41 2
474 184
442 184
1 0 15 0 0 4096 0 9 0 0 42 2
473 146
428 146
2 11 16 0 0 8320 0 8 1 0 0 4
474 239
364 239
364 74
338 74
2 13 17 0 0 4224 0 9 1 0 0 4
473 164
378 164
378 92
338 92
3 1 18 0 0 8320 0 15 4 0 0 4
523 117
543 117
543 146
549 146
1 0 19 0 0 4096 0 15 0 0 43 2
472 108
413 108
2 14 20 0 0 4224 0 15 1 0 0 4
472 126
384 126
384 101
338 101
3 0 21 0 0 8192 0 12 0 0 30 3
64 128
79 128
79 101
5 13 9 0 0 0 0 1 2 0 0 4
268 92
235 92
235 101
205 101
4 0 22 0 0 8320 0 10 0 0 37 3
254 225
217 225
217 47
0 2 23 0 0 4224 0 0 10 36 0 3
229 83
229 201
254 201
2 9 8 0 0 0 0 1 2 0 0 4
268 56
223 56
223 65
205 65
12 2 24 0 0 8320 0 1 7 0 0 4
338 83
371 83
371 202
474 202
6 0 21 0 0 0 0 2 0 0 30 2
141 101
133 101
3 3 21 0 0 12416 0 3 2 0 0 6
42 65
29 65
29 101
133 101
133 65
141 65
4 0 25 0 0 12416 0 3 0 0 32 4
42 74
37 74
37 92
118 92
5 8 25 0 0 0 0 2 3 0 0 4
141 92
118 92
118 74
112 74
4 7 26 0 0 8320 0 2 3 0 0 4
141 83
125 83
125 65
112 65
2 6 27 0 0 4224 0 2 3 0 0 2
141 56
112 56
1 5 28 0 0 4224 0 2 3 0 0 2
141 47
112 47
4 11 23 0 0 0 0 1 2 0 0 2
268 83
205 83
7 1 22 0 0 0 0 2 1 0 0 2
205 47
268 47
1 0 29 0 0 4096 0 16 0 0 39 2
457 306
457 318
1 1 29 0 0 8320 0 19 11 0 0 4
413 306
413 318
484 318
484 296
5 2 13 0 0 4224 0 14 16 0 0 2
457 94
457 270
2 8 14 0 0 4224 0 17 14 0 0 2
442 269
442 94
7 2 15 0 0 4224 0 14 18 0 0 2
428 94
428 269
6 2 19 0 0 4224 0 14 19 0 0 2
413 94
413 270
1 0 29 0 0 0 0 18 0 0 39 2
428 305
428 318
1 0 29 0 0 0 0 17 0 0 39 2
442 305
442 318
4 10 30 0 0 4224 0 14 1 0 0 2
384 65
338 65
3 9 15 0 0 12416 31 14 1 0 0 4
384 50
378 50
378 56
338 56
2 8 32 0 0 12416 0 14 1 0 0 4
384 36
372 36
372 47
338 47
7 1 33 0 0 4224 0 1 14 0 0 4
338 38
364 38
364 21
384 21
0
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
