CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 715 397
7 5.000 V
7 5.000 V
3 GND
500 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 715 397
12058632 0
0
0
0
0
0
0
11
5 SAVE-
218 260 85 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
22 *Combine
*TRAN -20 20
0
0
0
3

0 0 0 -1610612600
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 150 82 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
22 *Combine
*TRAN -20 20
0
0
0
3

0 0 0 -1610612600
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
7 Ground~
168 74 134 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -1610612600
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
2 +V
167 196 158 0 1 64
0 6
0
0 0 53600 -19276
3 -9V
-10 2 11 10
2 V1
-6 -8 8 0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -1610612600
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
2 +V
167 196 74 0 1 64
0 5
0
0 0 53600 0
3 +9V
-11 -14 10 -6
2 V2
-7 -24 7 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -1610612600
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
7 Ground~
168 260 266 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -1610612600
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
8 Op-Amp5~
219 196 113 0 5 64
0 7 4 5 6 3
8 Op-Amp5~
0 0 320 0
5 LM348
11 -16 46 -8
3 U1A
19 -26 40 -18
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 DIP14
64

0 3 2 4 11 1 3 2 4 11
1 5 6 4 11 7 10 9 4 11
8 12 13 4 11 14 894 6007 0 28460
25942 4399 4097 -8372 21327 168 168 24656 2 184
176 2 -8344 9963 1956 1034 75 -8226 21327 1
0 28460 25678 6055 4097 21327 -8293 -32025 6079 -8226
21327 75 1034 1956 0
88 0 0 0 4 1 0 0
1 U
9914 0 0
0
0
10 Capacitor~
219 105 107 0 2 64
0 2 4
10 Capacitor~
0 0 832 0
5 .01uF
-19 -18 16 -10
1 C
-3 -29 4 -21
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -1610612600
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
9 Resistor~
219 207 40 0 2 64
0 4 3
9 Resistor~
0 0 864 0
4 100k
-13 -12 15 -4
1 R
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612672
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 260 156 0 2 64
0 7 3
9 Resistor~
0 0 352 90
4 100k
6 -3 34 5
2 R2
13 -13 27 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612600
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 260 223 0 3 64
0 2 7 -1
9 Resistor~
0 0 352 90
3 27k
8 -2 29 6
2 R3
11 -12 25 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612684
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
10
5 0 3 0 0 4096 0 7 0 0 10 2
214 113
260 113
1 0 4 0 0 8320 0 9 0 0 7 3
189 40
150 40
150 107
1 3 5 0 0 4224 0 5 7 0 0 2
196 83
196 100
1 4 6 0 0 4224 0 4 7 0 0 2
196 143
196 126
1 0 7 0 0 12416 0 7 0 0 9 4
178 119
150 119
150 190
260 190
1 1 2 0 0 4224 0 8 3 0 0 3
96 107
74 107
74 128
2 2 4 0 0 0 0 7 8 0 0 2
178 107
114 107
1 1 2 0 0 0 0 11 6 0 0 2
260 241
260 260
1 2 7 0 0 0 0 10 11 0 0 2
260 174
260 205
2 2 3 0 0 8320 0 9 10 0 0 3
225 40
260 40
260 138
0
0
16 0 1
0
0
2 VD
0 2 0.01
0
0 0 0
0 0 1 2
0 0.01 0.0001 0.0001
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3540 8550976 100 100 0 0
77 66 677 276
0 397 715 738
675 66
77 66
677 67
677 276
0 0
4.98491e-315 0 5.39262e-315 1.6003e-314 4.98503e-315 4.98503e-315
12409 0
4 0.003 5
2
260 69
0 3 0 0 2	0 10 0 0
150 69
0 4 0 0 2	0 2 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
