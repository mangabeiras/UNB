CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 30 300 90 9
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
100 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 259
12058624 0
0
0
0
0
0
0
11
11 Signal Gen~
195 55 132 0 24 64
0 7 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1101004800 1094713344 0
0 953267991 953267991 990057071 1028443341
20
0 20 12 0 0 0.0001 0.0001 0.002 0.05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
5 12/0V
-18 -30 17 -22
2 V2
-8 -40 6 -32
0
0
44 %D %1 %2 DC 0 PULSE(12 0 0 100u 100u 2m 50m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
5 SAVE-
218 163 136 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
20 *Combine
*TRAN 0 12
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SAVE-
218 128 127 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
20 *Combine
*TRAN 0 12
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
4 .IC~
207 312 113 0 1 3
0 3
0
0 0 54080 0
2 0V
-7 -15 7 -7
4 CMD1
-14 -25 14 -17
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
3 CMD
6153 0 0
0
0
7 Ground~
168 238 213 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
2 +V
167 278 63 0 1 3
0 4
0
0 0 54112 0
3 12V
12 -2 33 6
2 V1
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
10 555 Timer~
219 238 127 0 8 17
0 2 7 6 4 5 3 3 4
10 555 Timer~
0 0 12992 0
5 UA555
-17 -23 18 -15
2 U1
-7 -33 7 -25
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 -33686019
88 0 496 0 1 1 0 0
1 U
9914 0 0
0
0
10 Capacitor~
219 355 172 0 2 5
0 2 3
10 Capacitor~
0 0 832 90
3 1uF
11 0 32 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 1 0 0
1 C
3747 0 0
0
0
10 Capacitor~
219 285 169 0 2 5
0 2 5
10 Capacitor~
0 0 832 90
5 0.1uF
11 0 46 8
2 C2
22 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 1 0 0
1 C
3549 0 0
0
0
9 Resistor~
219 151 166 0 3 5
0 2 6 -1
9 Resistor~
0 0 864 90
3 10k
7 0 28 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 355 106 0 4 5
0 3 4 0 1
9 Resistor~
0 0 864 90
3 27k
7 0 28 8
2 R2
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
9325 0 0
0
0
15
1 0 3 0 0 4096 0 4 0 0 3 2
312 125
312 136
7 0 3 0 0 4096 0 7 0 0 3 3
270 127
285 127
285 136
6 0 3 0 0 4224 0 7 0 0 4 2
270 136
355 136
1 2 3 0 0 0 0 11 8 0 0 2
355 124
355 163
1 0 2 0 0 4096 0 5 0 0 9 2
238 207
238 194
1 0 2 0 0 0 0 10 0 0 9 2
151 184
151 194
1 0 2 0 0 4096 0 9 0 0 9 2
285 178
285 194
1 0 2 0 0 8192 0 7 0 0 9 3
206 118
193 118
193 194
1 2 2 0 0 8320 0 8 1 0 0 5
355 181
355 194
118 194
118 137
86 137
2 0 4 0 0 8192 0 11 0 0 13 3
355 88
355 78
278 78
5 2 5 0 0 4224 0 7 9 0 0 3
270 145
285 145
285 160
0 4 4 0 0 4224 0 0 7 13 0 4
278 85
182 85
182 145
206 145
8 1 4 0 0 0 0 7 6 0 0 3
270 118
278 118
278 72
3 2 6 0 0 4224 0 7 10 0 0 3
206 136
151 136
151 148
1 2 7 0 0 4224 0 1 7 0 0 2
86 127
206 127
2
-16 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 50
1 20 251 73
5 24 245 62
50 Negative Edge Triggered 
555 Mono-stable Circuit
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 28
6 57 238 81
10 61 234 77
28 R2 and C1 control the delay.
33 .OPTIONS ITL4=100.0 TRTOL=3.000

16 0 0
0
0
3 Vin
-1.5 -0.7 0.02
3 Vcc
10 14 1
100 0 1 1e+006
0 0.05 0.0002 0.0002
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2556 8550464 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
5.08119e-315 0 5.39824e-315 1.5915e-314 5.08119e-315 5.08119e-315
16 0
4 0.01 10
1
332 136
0 3 0 0 1	0 3 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
