CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
245 80 857 348
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 0 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
2 2 0.500000 0.500000
245 357 857 634
42991616 0
0
0
0
0
0
0
18
13 Logic Switch~
5 147 153 0 2 11
0 15 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
34 0 0
2
36626.4 0
0
13 Logic Switch~
5 147 168 0 2 11
0 16 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6357 0 0
2
36626.4 1
0
13 Logic Switch~
5 147 183 0 2 11
0 17 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
319 0 0
2
36626.4 2
0
13 Logic Switch~
5 147 198 0 2 11
0 18 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3976 0 0
2
36626.4 3
0
14 Ascii Display~
172 440 166 0 42 43
0 9 8 7 6 5 4 3 2 0
64 17260 26979 27424 28526 8308 26725 8224 8224 16723
17225 18720 27493 31008 24948 8308 26725 27749 26228 11296
29800 25966 8308 31088 25888 28526 8308 26725 8299 25977
25199 24946 25646
0
0 0 20592 0
4 1MEG
-15 -42 13 -34
2 R5
-8 -52 6 -44
0
0
102 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
%DE %5 0 %V
%DF %6 0 %V
%DG %7 0 %V
%DH %8 0 %V
0
0
0
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
82 0 0 0 1 0 0 0
4 DISP
7634 0 0
2
36626.4 4
0
6 74LS85
106 264 156 0 14 29
0 11 12 13 14 15 16 17 18 19
20 21 22 10 23
0
0 0 12784 0
6 74LS85
-21 -51 21 -43
2 A6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 -33686019
65 0 0 512 1 1 0 0
1 U
523 0 0
2
36626.4 5
0
14 Logic Display~
6 315 126 0 1 3
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 R7
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
36626.4 6
0
14 Logic Display~
6 450 22 0 1 3
15 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 R8
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6901 0 0
2
36626.4 7
0
14 Logic Display~
6 431 36 0 1 3
13 12
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 R9
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
842 0 0
2
36626.4 8
0
14 Logic Display~
6 413 52 0 1 3
12 13
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 R10
13 -26 34 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
36626.4 9
0
14 Logic Display~
6 393 66 0 1 3
10 14
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 R11
13 -26 34 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
36626.4 10
0
12 Hex Display~
7 271 36 0 16 19
10 14 13 12 11 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
3 R12
-12 -52 9 -44
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4720 0 0
2
36626.4 11
0
9 Data Seq~
170 69 44 0 17 21
0 24 25 26 27 11 12 13 14 28
29 1 1 16 1 2 0 17
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
3 A13
-11 -54 10 -46
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
0
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
5551 0 0
2
36626.4 12
0
AAAAABACADAEAFAGAHAIAJAKALAMANAOAP
5 SCOPE
12 163 21 0 1 3
0 14
0
0 0 61680 0
3 TP1
-11 -4 10 4
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6986 0 0
2
36626.4 13
0
5 SCOPE
12 188 36 0 1 3
0 13
0
0 0 61680 0
3 TP2
-11 -4 10 4
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8745 0 0
2
36626.4 14
0
5 SCOPE
12 211 51 0 1 3
0 12
0
0 0 61680 0
3 TP3
-11 -4 10 4
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9592 0 0
2
36626.4 15
0
5 SCOPE
12 236 66 0 1 3
0 11
0
0 0 61680 0
3 TP4
-11 -4 10 4
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8748 0 0
2
36626.4 16
0
10 Ascii Key~
169 76 169 0 11 11
0 3 4 5 6 7 8 9 2 0
0 46
0
0 0 20528 0
0
0
0
0
0
0
0
0
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
3 KBD
7168 0 0
2
36626.4 17
0
43
8 -145589 2 0 0 4096 0 5 0 0 26 2
368 197
341 197
7 -3263 3 0 0 4224 0 5 0 0 26 2
374 189
341 189
6 -3262 4 0 0 4224 0 5 0 0 26 2
374 180
341 180
5 -3261 5 0 0 4224 0 5 0 0 26 2
374 171
341 171
4 -3260 6 0 0 4224 0 5 0 0 26 2
374 162
341 162
3 -3259 7 0 0 4224 0 5 0 0 26 2
374 153
341 153
2 -3258 8 0 0 4224 0 5 0 0 26 2
374 144
341 144
1 -3257 9 0 0 4224 0 5 0 0 26 2
374 135
341 135
13 1 10 0 0 8320 0 6 7 0 0 3
296 183
315 183
315 144
1 4 11 0 0 4160 0 17 0 0 43 2
236 78
236 101
1 3 12 0 0 4160 0 16 0 0 43 2
211 63
211 101
1 2 13 0 0 4288 0 15 0 0 43 2
188 48
188 101
1 1 14 0 0 4288 0 14 0 0 43 2
163 33
163 101
5 4 11 0 0 8192 0 13 0 0 43 3
101 53
139 53
139 101
6 3 12 0 0 8192 0 13 0 0 43 3
101 62
130 62
130 101
7 2 13 0 0 0 0 13 0 0 43 3
101 71
121 71
121 101
8 1 14 0 0 0 0 13 0 0 43 3
101 80
112 80
112 101
1 -3263 3 0 0 0 0 18 0 0 26 2
97 193
97 221
2 -3262 4 0 0 0 0 18 0 0 26 2
91 193
91 221
3 -3261 5 0 0 0 0 18 0 0 26 2
85 193
85 221
4 -3260 6 0 0 0 0 18 0 0 26 2
79 193
79 221
5 -3259 7 0 0 0 0 18 0 0 26 2
73 193
73 221
6 -3258 8 0 0 0 0 18 0 0 26 2
67 193
67 221
7 -3257 9 0 0 0 0 18 0 0 26 2
61 193
61 221
8 -145589 2 0 0 4224 0 18 0 0 26 2
55 193
55 221
-177604 0 1 0 0 4128 0 0 0 0 0 3
37 221
341 221
341 124
1 1 14 0 0 64 0 12 0 0 43 2
280 60
280 101
2 2 13 0 0 64 0 12 0 0 43 2
274 60
274 101
3 3 12 0 0 4160 0 12 0 0 43 2
268 60
268 101
4 4 11 0 0 64 0 12 0 0 43 2
262 60
262 101
1 4 11 0 0 64 0 6 0 0 43 3
232 129
221 129
221 101
2 3 12 0 0 64 0 6 0 0 43 3
232 138
210 138
210 101
3 2 13 0 0 64 0 6 0 0 43 3
232 147
199 147
199 101
4 1 14 0 0 64 0 6 0 0 43 3
232 156
188 156
188 101
5 1 15 0 0 4224 0 6 1 0 0 4
232 165
179 165
179 153
159 153
1 6 16 0 0 12416 0 2 6 0 0 4
159 168
170 168
170 174
232 174
7 1 17 0 0 4224 0 6 3 0 0 2
232 183
159 183
1 8 18 0 0 12416 0 4 6 0 0 4
159 198
174 198
174 192
232 192
1 4 11 0 0 4288 0 8 0 0 43 2
450 40
450 101
1 3 12 0 0 4288 0 9 0 0 43 2
431 54
431 101
1 2 13 0 0 64 0 10 0 0 43 2
413 70
413 101
1 1 14 0 0 64 0 11 0 0 43 2
393 84
393 101
-144844 0 1 0 0 4256 0 0 0 0 0 2
40 101
473 101
3
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 10
59 100 175 124
63 104 157 128
10 Data Bus 1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
42 124 112 144
46 128 109 142
9 ASCII Key
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 10
181 201 246 222
185 205 243 220
10 Data Bus 2
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 100 100 0 0
77 66 977 246
0 0 0 0
977 66
77 66
977 66
977 246
0 0
4.94359e-315 0 5.30706e-315 1.5917e-314 4.94359e-315 4.94359e-315
12401 0
0 0.001 2
0
0 0 100 100 0 0
77 66 977 246
0 0 0 0
977 66
77 66
977 66
977 246
0 0
4.94359e-315 0 5.30499e-315 1.58735e-314 4.94359e-315 4.94359e-315
12401 0
0 0.001 0.5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
