CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
15 0 15 100 3
25 103 545 447
7 5.000 V
7 5.000 V
3 GND
25 103 545 447
142606338 0
0
0
0
0
0
0
5
13 Logic Switch~
5 61 250 0 2 3
0 2 -99
0
0 0 20576 0
2 0V
-7 -16 7 -8
2 S1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 62 156 0 2 3
0 3 -99
0
0 0 20576 0
2 0V
-7 -16 7 -8
2 S2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
13 Piezo Buzzer~
174 106 203 0 2 5
10 3 2
0
0 0 4192 270
4 .1uF
10 -16 38 -8
3 BZ1
13 -26 34 -18
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
2 BZ
3618 0 0
0
0
9 Data Seq~
170 67 67 0 17 21
0 6 7 8 9 10 11 4 5 12
13 3 1 4 25 16 0 33
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -54 10 -46
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
0
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 0 0 0 0
2 DS
6153 0 0
0
0
AAAAABAAACAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
8 Speaker~
175 196 68 0 2 5
10 4 5
0
0 0 20576 0
1 8
-3 -22 4 -14
0
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
3 SPK
5394 0 0
0
0
4
1 2 2 0 0 4224 0 1 3 0 0 3
73 250
106 250
106 234
1 1 3 0 0 4224 0 2 3 0 0 3
74 156
106 156
106 172
1 7 4 0 0 12416 0 5 4 0 0 5
188 52
188 39
137 39
137 94
99 94
8 2 5 0 0 4224 0 4 5 0 0 3
99 103
188 103
188 84
0
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
