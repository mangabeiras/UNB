CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 594 357
7 5.000 V
7 5.000 V
3 GND
0 66 594 357
12058626 0
0
0
0
0
0
0
12
5 SAVE-
218 219 60 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 C
3 -26 10 -18
0
0
0
24 *Combine
*TRAN -170 500
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
11 Signal Gen~
195 64 123 0 24 64
0 6 2 5 86 -8 8 5 0 0
0 0 0 0 0 0 0 994360628 0 0
994352038 0 994356333 1133903872 994360628
20
0 0.003002 0 0 0.003 0 0.003001 300 0.003002 0
0 0 0 0 0 0 0 0 0 0
0
0 0 16704 0
6 0/300V
-20 -28 22 -20
2 V1
-6 -38 8 -30
0
0
48 %D %1 %2 DC 0 PWL( 0 0 3m 0 3.001m 300 3.002m 0)
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
5 SAVE-
218 119 175 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
10 *TRAN -1 6
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
11 Signal Gen~
195 64 180 0 24 64
0 8 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1123031187 0 1084227584
1002740646 869711765 869711765 981668463 1007188621
20
0 120.048 0 5 0.006 1e-007 1e-007 0.001 0.00833 0
0 0 0 0 0 0 0 0 0 0
0
0 0 16704 0
4 0/5V
-14 -28 14 -20
2 V2
-7 -38 7 -30
0
0
46 %D %1 %2 DC 0 PULSE(0 5 6m 100n 100n 1m 8.33m)
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
5 SAVE-
218 234 136 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
24 *Combine
*TRAN -170 500
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
7 Ground~
168 106 208 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
11 Signal Gen~
195 64 65 0 19 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1114636288 0 1126825984
20
1 60 0 170 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 16704 0
9 -170/170V
-30 -28 33 -20
2 V3
-7 -38 7 -30
0
0
38 %D %1 %2 DC 0 SIN(0 170 60 0 0) AC 1 0
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
7 Ground~
168 233 207 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
8 V-Math2~
219 165 69 0 3 64
0 7 6 5
8 V-Math2~
0 0 5184 0
4 ADDV
-14 -36 14 -27
2 M1
-7 -46 7 -38
6 V(A+B)
-21 -24 21 -16
0
14 %D %1 %2 %3 %S
0
0
6 V(A+B)
7

0 1 2 3 1 2 3 -33686019
88 0 0 0 1 0 0 0
1 M
3549 0 0
0
0
8 Triac:B~
219 233 165 0 3 64
0 4 3 2
8 Triac:B~
0 0 320 0
8 MAC210-6
20 -4 76 4
2 Q1
41 -14 55 -6
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-220
7

0 2 3 1 2 3 1 -33686019
88 0 0 0 1 0 0 0
1 Q
7931 0 0
0
0
9 Resistor~
219 160 175 0 2 64
0 8 3
9 Resistor~
0 0 352 0
2 50
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 233 91 0 2 64
0 5 4
9 Resistor~
0 0 352 270
3 100
5 -2 26 6
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
10
3 1 2 0 0 4096 0 10 8 0 0 2
233 183
233 201
2 2 3 0 0 4224 0 10 11 0 0 2
217 175
178 175
2 1 4 0 0 4224 0 12 10 0 0 2
233 109
233 147
1 3 5 0 0 8320 0 12 9 0 0 3
233 73
233 60
199 60
1 2 6 0 0 8320 0 2 9 0 0 4
95 118
123 118
123 69
131 69
2 0 2 0 0 0 0 2 0 0 8 2
95 128
106 128
2 0 2 0 0 0 0 4 0 0 8 2
95 185
106 185
2 1 2 0 0 8320 0 7 6 0 0 3
95 70
106 70
106 202
1 1 7 0 0 4224 0 9 7 0 0 2
131 60
95 60
1 1 8 0 0 4224 0 4 11 0 0 2
95 175
142 175
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 214
286 4 550 148
290 8 546 120
214 In this circuit, a piecewise 
generator creates an 
"industrial spike" which is 
then added to the AC source. 
This spike causes the triac to 
fire prematurely (before it is 
gated on by the 5V pulser).
0
17 0 1
0
0
2 IA
-0.02 0.02 0.0001
0
0 0 0
0 0 1 2
0 0.04333 0.0004167 0.0004167 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
