CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 100 3
0 66 640 343
7 5.000 V
7 5.000 V
3 GND
0 343 640 452
159383554 0
0
0
0
0
0
0
9
13 Logic Switch~
5 55 130 0 2 3
0 2 -99
0
0 0 20576 0
2 0V
-7 -16 7 -8
2 S1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 56 106 0 2 3
0 6 -99
0
0 0 20576 0
2 0V
-7 -16 7 -8
2 S2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
11 SPDT Relay~
176 113 111 0 10 11
0 5 4 3 6 2 0 0 0 0
1
0
0 0 20832 0
7 12VSPDT
-27 -35 22 -27
4 RLY1
21 -2 49 6
0
0
20 %D %1 %2 %3 %4 %5 %S
0
45 alias:XSPDTRELAY {PULLIN=9.6 RESISTANCE=1000}
4 DIP4
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 0 0 0 0 0
3 RLY
3618 0 0
0
0
14 Logic Display~
6 209 37 0 1 3
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 150 38 0 1 3
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
5 SCOPE
12 342 64 0 3 3
0 2 99 49
0
0 0 57568 0
1 1
-4 -4 3 4
2 V1
-7 -14 7 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 300 64 0 3 3
0 3 99 50
0
0 0 57568 0
1 2
-4 -4 3 4
2 V2
-7 -14 7 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 257 64 0 3 3
0 4 99 51
0
0 0 57568 0
1 3
-4 -4 3 4
2 V3
-7 -14 7 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3747 0 0
0
0
2 +V
167 178 53 0 1 3
0 5
0
0 0 53728 0
3 10V
-11 -22 10 -14
2 V4
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3549 0 0
0
0
8
0 1 2 0 0 8320 0 0 6 7 0 4
90 130
90 147
342 147
342 76
1 0 3 0 0 4096 0 4 0 0 5 2
209 55
209 100
1 0 4 0 0 4096 0 5 0 0 6 2
150 56
150 86
1 1 5 0 0 4224 0 3 9 0 0 3
127 93
178 93
178 62
1 3 3 0 0 8320 0 7 3 0 0 3
300 76
300 100
127 100
2 1 4 0 0 4224 0 3 8 0 0 3
127 86
257 86
257 76
5 1 2 0 0 0 0 3 1 0 0 2
97 130
67 130
4 1 6 0 0 4224 0 3 2 0 0 2
97 106
68 106
0
0
16 2 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.001 5e-005 5e-005 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
1348 8550464 100 100 0 0
77 66 287 216
320 66 640 354
286 66
77 66
287 66
287 216
0 0
4.85009e-315 0 4.85857e-315 0 4.85009e-315 4.85857e-315
16 0
4 0.0003 5
1
209 74
0 3 0 0 1	0 2 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
