CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 373 402
7 5.000 V
7 5.000 V
3 GND
2500 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 373 402
9961472 0
0
0
0
0
0
0
19
5 SAVE-
218 192 87 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
24 *Combine
*DC -614m 11.9
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 145 87 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
24 *Combine
*DC -614m 11.9
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
7 Ground~
168 77 155 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
11 Signal Gen~
195 36 114 0 19 64
0 9 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1036831949
20
1 1000 0 0.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 576 0
11 -100m/100mV
-36 -48 41 -40
3 Vin
-14 -35 7 -27
0
0
39 %D %1 %2 DC 0 SIN(0 100m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
7 Ground~
168 284 212 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
2 +V
167 169 274 0 1 64
0 3
0
0 0 54112 180
4 -12V
3 4 31 12
3 Vee
-24 3 -3 11
0
4 Vee;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
2 +V
167 170 19 0 1 64
0 4
0
0 0 54112 0
3 12v
6 -14 27 -6
3 Vcc
-18 -13 3 -5
0
4 VCC;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
10 NPN Trans~
219 138 109 0 3 64
0 13 14 11
10 NPN Trans~
0 0 832 0
7 2N2222A
-46 14 3 22
2 Q1
-21 3 -7 11
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 -33686019
81 0 0 0 1 1 0 0
1 Q
3747 0 0
0
0
10 NPN Trans~
219 199 110 0 3 64
0 5 12 11
10 NPN Trans~
0 0 832 512
7 2N2222A
1 12 50 20
2 Q2
9 2 23 10
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 -33686019
81 0 0 0 1 1 0 0
1 Q
3549 0 0
0
0
10 NPN Trans~
219 176 173 0 3 64
0 11 6 10
10 NPN Trans~
0 0 832 512
7 2N2222A
-56 -1 -7 7
2 Q3
-38 -11 -24 -3
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 -33686019
81 0 0 0 1 1 0 0
1 Q
7931 0 0
0
0
6 Diode~
219 228 195 0 2 64
0 6 7
6 Diode~
0 0 832 270
5 1N914
9 0 44 8
2 D1
18 -10 32 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
9325 0 0
0
0
6 Diode~
219 228 227 0 2 64
0 7 8
6 Diode~
0 0 832 270
5 1N914
13 2 48 10
2 D2
21 -7 35 1
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
8903 0 0
0
0
9 Resistor~
219 145 63 0 4 64
0 13 4 0 1
9 Resistor~
0 0 4960 90
5 7.75k
-41 6 -6 14
3 RC1
-33 -6 -12 2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 192 63 0 4 64
0 5 4 0 1
9 Resistor~
0 0 4960 602
5 7.75k
7 0 42 8
3 RC2
14 -10 35 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 252 110 0 4 64
0 12 2 0 -1
9 Resistor~
0 0 4960 0
2 50
-7 -12 7 -4
3 RB2
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 96 109 0 2 64
0 9 14
9 Resistor~
0 0 4960 0
2 50
-7 -12 7 -4
3 RB1
-10 -23 11 -15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 169 217 0 3 64
0 3 10 1
9 Resistor~
0 0 4960 90
4 2.5k
-32 0 -4 8
2 RE
-25 -10 -11 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 200 247 0 4 64
0 8 3 0 1
9 Resistor~
0 0 4960 180
4 1.5k
-14 -12 14 -4
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 256 173 0 4 64
0 6 2 0 -1
9 Resistor~
0 0 4960 0
4 3.2k
-14 -12 14 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
19
1 1 5 0 0 4224 0 9 14 0 0 2
192 92
192 81
2 1 2 0 0 8192 0 4 3 0 0 3
67 119
77 119
77 149
1 0 6 0 0 4096 0 11 0 0 6 2
228 185
228 173
2 0 2 0 0 0 0 19 0 0 5 2
274 173
284 173
2 1 2 0 0 8320 0 15 5 0 0 3
270 110
284 110
284 206
2 1 6 0 0 4224 0 10 19 0 0 2
182 173
238 173
1 2 7 0 0 4224 0 12 11 0 0 2
228 217
228 205
2 1 8 0 0 4224 0 12 18 0 0 3
228 237
228 247
218 247
0 2 3 0 0 4096 0 0 18 11 0 2
169 247
182 247
1 1 9 0 0 4224 0 16 4 0 0 4
78 109
63 109
63 109
67 109
1 1 3 0 0 4224 0 17 6 0 0 2
169 235
169 259
3 2 10 0 0 4224 0 10 17 0 0 2
169 191
169 199
1 0 11 0 0 4096 0 10 0 0 14 2
169 155
169 139
3 3 11 0 0 8320 0 9 8 0 0 4
192 128
192 139
145 139
145 127
2 1 12 0 0 4224 0 9 15 0 0 2
205 110
234 110
1 0 4 0 0 4096 0 7 0 0 17 2
170 28
170 36
2 2 4 0 0 8320 0 13 14 0 0 4
145 45
145 36
192 36
192 45
1 1 13 0 0 4224 0 8 13 0 0 2
145 91
145 81
2 2 14 0 0 4224 0 16 8 0 0 2
114 109
132 109
0
21 .OPTIONS METHOD=GEAR

4 0 0
0
0
3 Vin
-0.1 0.1 0.01
3 Vee
-15 0 1
100 0 1 1e+006
0 0.002 2.5e-005 2.5e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
