CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 27 100 9
0 66 548 396
7 5.000 V
7 5.000 V
3 GND
5e+006 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 548 396
11010066 1
0
0
0
0
0
0
6
7 Ground~
168 241 191 0 64 64
0 2 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
11 Multimeter~
205 119 64 0 64 64
0 2 6 7 5 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
4 73 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
0
0 0 16448 0
6 1.000u
-21 -19 21 -11
4 I0m1
-14 -29 14 -21
0
0
31 R1%D %1 %2 1E-9
%D %4 %2 DC %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
73 0 0 0 1 1 0 0
1 I
4441 0 0
0
0
9 Resistor~
219 271 92 0 64 64
0 4 3 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
9 Resistor~
0 0 352 0
2 1k
-7 -12 7 -4
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
9 Resistor~
219 191 92 0 64 64
0 5 4 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
9 Resistor~
0 0 352 0
3 500
-10 -12 11 -4
2 R3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
9 Resistor~
219 354 92 0 64 64
0 3 2 0 -1 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
9 Resistor~
0 0 352 0
2 2K
-7 -12 7 -4
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 273 123 0 64 64
0 4 3 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
9 Resistor~
0 0 352 0
2 1k
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
7
1 0 2 0 0 4096 0 1 0 0 2 2
241 185
241 172
2 1 2 0 0 12416 0 5 2 0 0 5
372 92
387 92
387 172
94 172
94 87
2 0 3 0 0 8192 0 6 0 0 4 3
291 123
316 123
316 92
2 1 3 0 0 4224 0 3 5 0 0 2
289 92
336 92
1 0 4 0 0 8192 0 6 0 0 6 3
255 123
233 123
233 92
2 1 4 0 0 4224 0 4 3 0 0 2
209 92
253 92
4 1 5 0 0 8320 0 2 4 0 0 3
144 87
144 92
173 92
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-006 1e-007 1e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1292 1210432 100 100 0 0
0 0 0 0
7 90 147 160
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
4 0.001 0.002
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
