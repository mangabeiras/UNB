CircuitMaker Text
5.5
41 91 70 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 27 100 9
12 70 613 451
8  5.000 V
8  5.000 V
3 GND
1000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
12 70 613 451
8388626 0
0
0
0
0
0
0
20
13 Logic Switch~
5 65 278 0 1 11
0 13
0
0 0 4448 0
2 5V
-7 -16 7 -8
2 S1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 64 157 0 1 11
0 16
0
0 0 4448 0
2 5V
-7 -16 7 -8
2 S2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 63 108 0 1 11
0 17
0
0 0 4448 0
2 5V
-7 -16 7 -8
2 S3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
10 3-In NAND~
219 324 300 0 4 21
0 13 12 11 3
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U2A
-13 -4 8 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 -33686019
65 0 0 0 3 1 6 0
1 U
6153 0 0
0
0
10 3-In NAND~
219 324 247 0 4 21
0 14 12 13 4
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U3C
-13 -4 8 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 -33686019
65 0 0 0 3 3 7 0
1 U
5394 0 0
0
0
10 3-In NAND~
219 322 181 0 4 21
0 15 11 13 5
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U3B
-12 -4 9 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 -33686019
65 0 0 0 3 2 7 0
1 U
7734 0 0
0
0
10 3-In NAND~
219 321 117 0 4 21
0 15 14 13 6
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U3A
-13 -3 8 5
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 -33686019
65 0 0 0 3 1 7 0
1 U
9914 0 0
0
0
9 Inverter~
13 221 157 0 2 21
0 11 14
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1D
-7 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 4 5 0
1 U
3747 0 0
0
0
9 Inverter~
13 220 108 0 2 21
0 12 15
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1C
-8 -22 13 -14
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 3 5 0
1 U
3549 0 0
0
0
9 Inverter~
13 122 157 0 2 21
0 16 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1B
-7 -22 14 -14
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 2 5 0
1 U
7931 0 0
0
0
9 Inverter~
13 121 108 0 2 21
0 17 12
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1A
-7 -22 14 -14
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 1 5 0
1 U
9325 0 0
0
0
2 +V
167 465 17 0 1 3
0 2
0
0 0 53472 0
3 10V
12 -2 33 6
2 V1
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
4 LED~
171 537 105 0 2 5
10 7 3
0
0 0 96 0
4 LED2
10 -16 38 -8
2 D1
17 -26 31 -18
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3834 0 0
0
0
4 LED~
171 488 106 0 2 5
10 8 4
0
0 0 96 0
4 LED2
10 -16 38 -8
2 D2
17 -26 31 -18
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3363 0 0
0
0
4 LED~
171 435 107 0 2 5
10 9 5
0
0 0 96 0
4 LED2
10 -16 38 -8
2 D3
17 -26 31 -18
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7668 0 0
0
0
4 LED~
171 382 106 0 2 5
10 10 6
0
0 0 96 0
4 LED2
10 -16 38 -8
2 D4
17 -26 31 -18
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4718 0 0
0
0
9 Resistor~
219 382 66 0 4 5
0 10 2 0 1
9 Resistor~
0 0 96 90
2 1k
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 435 66 0 4 5
0 9 2 0 1
9 Resistor~
0 0 96 90
2 1k
-7 -12 7 -4
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 488 67 0 4 5
0 8 2 0 1
9 Resistor~
0 0 96 90
2 1k
-7 -12 7 -4
2 R3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 537 67 0 4 5
0 7 2 0 1
9 Resistor~
0 0 96 90
2 1k
-7 -12 7 -4
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
4871 0 0
0
0
28
1 0 2 0 0 4096 0 12 0 0 4 2
465 26
465 35
2 0 2 0 0 4096 0 18 0 0 4 2
435 48
435 35
2 0 2 0 0 4096 0 19 0 0 4 2
488 49
488 35
2 2 2 0 0 8320 0 17 20 0 0 4
382 48
382 35
537 35
537 49
2 4 3 0 0 8320 0 13 4 0 0 3
537 115
537 300
351 300
2 4 4 0 0 8320 0 14 5 0 0 3
488 116
488 247
351 247
2 4 5 0 0 8320 0 15 6 0 0 3
435 117
435 181
349 181
2 4 6 0 0 8320 0 16 7 0 0 3
382 116
382 117
348 117
1 1 7 0 0 4224 0 20 13 0 0 2
537 85
537 95
1 1 8 0 0 4224 0 19 14 0 0 2
488 85
488 96
1 1 9 0 0 4224 0 18 15 0 0 2
435 84
435 97
1 1 10 0 0 4224 0 17 16 0 0 2
382 84
382 96
2 0 11 0 0 4096 0 6 0 0 16 2
298 181
171 181
2 0 12 0 0 4096 0 5 0 0 17 2
300 247
181 247
1 0 13 0 0 4224 0 1 0 0 20 2
77 278
275 278
0 3 11 0 0 4224 0 0 4 25 0 3
171 157
171 309
300 309
0 2 12 0 0 4224 0 0 4 26 0 3
181 108
181 300
300 300
3 0 13 0 0 0 0 5 0 0 20 2
300 256
275 256
3 0 13 0 0 0 0 6 0 0 20 2
298 190
275 190
3 1 13 0 0 0 0 7 4 0 0 4
297 126
275 126
275 291
300 291
2 0 14 0 0 4096 0 8 0 0 22 2
242 157
283 157
2 1 14 0 0 8320 0 7 5 0 0 4
297 117
283 117
283 238
300 238
0 1 15 0 0 4224 0 0 6 24 0 3
267 108
267 172
298 172
2 1 15 0 0 0 0 9 7 0 0 2
241 108
297 108
2 1 11 0 0 0 0 10 8 0 0 2
143 157
206 157
2 1 12 0 0 0 0 11 9 0 0 2
142 108
205 108
1 1 16 0 0 4224 0 2 10 0 0 2
76 157
107 157
1 1 17 0 0 4224 0 3 11 0 0 2
75 108
106 108
0
31 .OPTIONS METHOD=GEAR MAXORD=2

2049 0 0
0
0
3 Vin
-0.1 0.1 0.005
3 Vee
-15 0 1
100 0 1 1e+006
0 0.005 2.5e-005 2.5e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1324 1210432 100 100 0 0
0 0 0 0
1 57 141 127
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
16 0
4 2 2
1
406 300
0 4 0 0 2	0 5 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
