CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 325
7 5.000 V
7 5.000 V
3 GND
0 66 640 325
9961474 0
0
0
0
0
0
0
21
7 Ground~
168 111 138 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
7 Trans3~
219 161 104 0 5 11
0 11 2 5 2 4
0
0 0 336 0
6 5TO1CT
-20 -32 22 -24
2 T1
-6 -42 8 -34
0
0
20 %D %1 %2 %3 %4 %5 %S
0
25 alias:XTRANSCT {RATIO=.2}
0
11

0 1 2 3 4 5 1 2 3 4
5 0
88 0 0 0 1 0 0 0
1 T
4441 0 0
0
0
5 SAVE-
218 545 179 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 D
3 -26 10 -18
0
0
0
21 *Combine
*TRAN -17 0
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SAVE-
218 540 27 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 C
3 -26 10 -18
0
0
0
20 *Combine
*TRAN 0 17
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
5 SAVE-
218 350 179 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
21 *Combine
*TRAN -17 0
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SAVE-
218 349 27 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
20 *Combine
*TRAN 0 17
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
10 Polar Cap~
219 525 60 0 2 5
0 6 2
10 Polar Cap~
0 0 848 26894
5 100uF
10 4 45 12
2 C1
21 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
9914 0 0
0
0
10 Polar Cap~
219 340 137 0 2 5
0 2 9
10 Polar Cap~
0 0 848 270
5 100uF
10 4 45 12
2 C2
21 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
3747 0 0
0
0
12 Zener Diode~
219 461 127 0 2 5
0 7 2
12 Zener Diode~
0 0 848 90
6 1N4736
14 -2 56 6
2 D1
28 -12 42 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
100 0 0 0 1 1 0 0
1 D
3549 0 0
0
0
10 Polar Cap~
219 340 57 0 2 5
0 10 2
10 Polar Cap~
0 0 848 270
5 100uF
10 4 45 12
2 C3
21 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
7931 0 0
0
0
12 Zener Diode~
219 461 82 0 2 5
0 2 8
12 Zener Diode~
0 0 848 90
6 1N4736
14 -2 56 6
2 D2
28 -12 42 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
100 0 0 0 1 1 0 0
1 D
9325 0 0
0
0
7 Ground~
168 595 120 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
10 FW Bridge~
219 258 89 0 4 9
0 9 5 10 4
10 FW Bridge~
0 0 848 90
6 BRIDGE
12 -34 54 -26
2 D3
21 -44 35 -36
0
0
17 %D %1 %2 %3 %4 %S
0
0
0
9

0 1 2 3 4 1 2 3 4 0
88 0 0 256 1 0 0 0
1 D
3834 0 0
0
0
11 Signal Gen~
195 40 98 0 19 64
0 11 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1114636288 0 1126825984
20
1 60 0 170 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 16976 0
9 -170/170V
-31 -28 32 -20
2 V1
-7 -38 7 -30
0
0
38 %D %1 %2 DC 0 SIN(0 170 60 0 0) AC 1 0
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
12 NPN Trans:C~
219 465 34 0 3 7
0 10 8 6
12 NPN Trans:C~
0 0 848 90
6 2N3904
-31 -27 11 -19
2 Q1
-31 -17 -17 -9
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
7668 0 0
0
0
12 PNP Trans:C~
219 465 172 0 3 7
0 9 7 3
12 PNP Trans:C~
0 0 848 27406
6 2N3906
-23 30 19 38
2 Q2
-9 20 5 28
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
113 0 0 0 1 1 0 0
1 Q
4718 0 0
0
0
10 Polar Cap~
219 525 149 0 2 5
0 2 3
10 Polar Cap~
0 0 848 26894
5 100uF
10 4 45 12
2 C4
21 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
3874 0 0
0
0
9 Resistor~
219 574 156 0 4 5
0 3 2 0 -1
9 Resistor~
0 0 4976 90
3 500
7 0 28 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 423 145 0 2 5
0 9 7
9 Resistor~
0 0 4976 0
3 680
-10 -12 11 -4
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 574 63 0 3 5
0 2 6 -1
9 Resistor~
0 0 4976 90
3 500
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 427 60 0 2 5
0 8 10
9 Resistor~
0 0 4976 180
3 680
-10 -12 11 -4
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3750 0 0
0
0
28
1 0 2 0 0 4096 0 1 0 0 20 2
111 132
111 115
3 1 3 0 0 4224 0 16 18 0 0 3
481 179
574 179
574 174
4 5 4 0 0 12416 0 13 2 0 0 4
292 85
299 85
299 123
183 123
2 3 5 0 0 4224 0 13 2 0 0 2
228 85
183 85
1 0 6 0 0 4096 0 7 0 0 19 2
524 50
524 27
0 2 2 0 0 4096 0 0 7 22 0 2
524 102
524 67
2 0 3 0 0 0 0 17 0 0 2 2
524 156
524 179
1 0 2 0 0 4096 0 17 0 0 22 2
524 139
524 102
2 0 2 0 0 0 0 9 0 0 22 2
463 115
463 102
1 0 2 0 0 0 0 11 0 0 22 2
463 90
463 102
1 0 2 0 0 0 0 20 0 0 22 2
574 81
574 102
2 0 2 0 0 0 0 18 0 0 22 2
574 138
574 102
2 0 7 0 0 4224 0 19 0 0 16 2
441 145
463 145
1 0 8 0 0 4096 0 21 0 0 15 2
445 60
463 60
2 2 8 0 0 4224 0 11 15 0 0 2
463 70
463 50
2 1 7 0 0 0 0 16 9 0 0 2
463 156
463 135
0 1 9 0 0 4096 0 0 19 24 0 3
395 179
395 145
405 145
0 2 10 0 0 4096 0 0 21 26 0 3
395 27
395 60
409 60
3 2 6 0 0 4224 0 15 20 0 0 3
481 27
574 27
574 45
2 2 2 0 0 4096 0 2 14 0 0 4
143 115
86 115
86 103
71 103
0 4 2 0 0 12288 0 0 2 22 0 6
339 102
312 102
312 160
216 160
216 104
183 104
1 0 2 0 0 8320 0 12 0 0 27 3
595 114
595 102
339 102
2 0 9 0 0 4096 0 8 0 0 24 2
339 144
339 179
1 1 9 0 0 8320 0 13 16 0 0 3
260 117
260 179
445 179
1 0 10 0 0 0 0 10 0 0 26 2
339 47
339 27
3 1 10 0 0 8320 0 13 15 0 0 3
260 53
260 27
445 27
2 1 2 0 0 0 0 10 8 0 0 2
339 64
339 127
1 1 11 0 0 4224 0 14 2 0 0 2
71 93
143 93
1
-16 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 22
2 5 232 34
7 9 227 28
22 +/-6 Volt Power Supply
23 .OPTIONS ABSTOL=1.000u

16 0 0
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 0.08333 0.0004167 0.0004167 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
3344 8526400 100 100 0 0
98 66 608 126
0 259 640 452
608 66
98 66
608 66
608 126
0 0
0.08333 0 18 -18 0.08333 0.08333
12409 0
4 0.02 100
5
518 27
0 6 0 0 1	0 19 0 0
514 179
0 3 0 0 1	0 2 0 0
369 27
0 10 0 0 2	0 26 0 0
204 85
0 5 0 0 1	0 4 0 0
372 179
0 9 0 0 2	0 24 0 0
0 0 100 100 0 0
77 66 617 126
0 0 0 0
617 66
77 66
617 66
617 126
0 0
0.0003 0 5 0 0.0003 0.0003
13433 0
0 5e-005 5
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
-0.72 -1.5 12.6 7.2 0.78 0.78
0 0
0 0.3 1e+036
0
0 0 100 100 0 0
77 66 293 126
0 0 0 0
293 66
77 66
293 66
293 126
0 0
1e+006 1 -3.55271e-015 -3.55271e-015 999999 999999
4211 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
