CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
100000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 259
9961474 0
0
0
0
0
0
0
14
7 Ground~
168 438 171 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
5 SAVE-
218 84 110 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
22 *Combine
*TRAN -30 20
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SAVE-
218 366 152 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
22 *Combine
*TRAN -30 20
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
7 Ground~
168 110 169 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
11 Signal Gen~
195 41 115 0 24 64
0 4 2 1 86 -7 7 0 0 0
0 0 0 0 0 0 0 1232348160 0 1097859072
0 869711765 869711765 886488981 897988541
20
0 1e+006 0 15 0 1e-007 1e-007 4e-007 1e-006 0
0 0 0 0 0 0 0 0 0 0
0
0 0 320 0
5 0/15V
-17 -28 18 -20
2 V1
-7 -38 7 -30
0
0
45 %D %1 %2 DC 0 PULSE(0 15 0 100n 100n 400n 1u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
6 Diode~
219 294 117 0 2 5
0 5 6
6 Diode~
0 0 64 26894
5 DIODE
-17 -18 18 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
7734 0 0
0
0
6 Diode~
219 355 119 0 2 5
0 3 5
6 Diode~
0 0 64 90
5 DIODE
-17 -18 18 -10
2 D2
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
9914 0 0
0
0
10 Capacitor~
219 268 84 0 2 5
0 7 5
10 Capacitor~
0 0 320 0
3 1uF
-12 -18 9 -10
2 C1
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
3747 0 0
0
0
10 Capacitor~
219 325 152 0 2 5
0 6 3
10 Capacitor~
0 0 320 0
3 1uF
-12 -18 9 -10
2 C2
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
3549 0 0
0
0
6 Diode~
219 172 117 0 2 5
0 7 2
6 Diode~
0 0 64 26894
5 DIODE
-17 -18 18 -10
2 D3
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
7931 0 0
0
0
6 Diode~
219 233 120 0 2 5
0 6 7
6 Diode~
0 0 64 90
5 DIODE
-17 -18 18 -10
2 D4
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
9325 0 0
0
0
10 Capacitor~
219 145 84 0 2 5
0 4 7
10 Capacitor~
0 0 320 0
3 1uF
-12 -18 9 -10
2 C3
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
8903 0 0
0
0
10 Capacitor~
219 203 152 0 2 5
0 2 6
10 Capacitor~
0 0 320 0
3 1uF
-12 -18 9 -10
2 C4
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
3834 0 0
0
0
9 Resistor~
219 408 152 0 4 5
0 3 2 0 -1
9 Resistor~
0 0 352 0
4 1Meg
-14 -12 14 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3363 0 0
0
0
15
2 0 2 0 0 4096 0 10 0 0 2 2
172 127
172 152
1 0 2 0 0 4224 0 13 0 0 6 2
194 152
110 152
1 0 3 0 0 4096 0 7 0 0 4 2
355 129
355 152
2 1 3 0 0 4224 0 9 14 0 0 2
334 152
390 152
2 1 2 0 0 0 0 14 1 0 0 3
426 152
438 152
438 165
2 1 2 0 0 0 0 5 4 0 0 3
72 120
110 120
110 163
1 1 4 0 0 12416 0 12 5 0 0 4
136 84
110 84
110 110
72 110
1 0 5 0 0 4096 0 6 0 0 13 2
294 107
294 84
2 0 6 0 0 4096 0 6 0 0 15 2
294 127
294 152
1 0 6 0 0 0 0 11 0 0 15 2
233 130
233 152
2 0 7 0 0 4096 0 11 0 0 14 2
233 110
233 84
1 0 7 0 0 0 0 10 0 0 14 2
172 107
172 84
2 2 5 0 0 4224 0 8 7 0 0 3
277 84
355 84
355 109
2 1 7 0 0 4224 0 12 8 0 0 2
154 84
259 84
2 1 6 0 0 4224 0 13 9 0 0 2
212 152
316 152
2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 168
18 190 354 274
22 194 350 258
168 The rail voltage (15V) is multiplied by 
each set of 2 diodes and 2 capacitors.  
Two sets have been used in this circuit 
resulting in a -30VDC (approx.) output.
-16 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 18
17 8 207 37
21 12 201 31
18 Voltage Multiplier
22 .OPTIONS BOOLH=15.00

17 0 1
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 5e-005 2.5e-008 2.5e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3456 1210432 100 100 0 0
98 66 608 126
323 79 463 149
608 66
77 66
617 66
617 126
0 0
0 0 0 0 0 0
16 0
4 1 2e-019
1
374 152
0 3 0 0 1	0 4 0 0
2500 8550464 100 100 0 0
77 66 617 126
-2 261 638 454
617 66
77 66
617 66
617 126
0 0
0 0 0 0 0 0
16 0
4 1e-005 100
1
385 152
0 3 0 0 1	0 4 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
