CircuitMaker Text
4
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 1e+012
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 0
0 66 624 296
0 66 624 296
144179202 2
0
0
0
0
0
0
15
5 SAVE-
218 493 106 0 11 
0 0 0 0 0 0 0 0 0 0 
1 0 0
0 0 -8000 0
1 D
3 -26 10 -18
0
0
0
20 *Combine
*TRAN 5u 5
0
1

0 0 
0 0 0 0 0 0 0 0
0
8953 0 0 0
5 SAVE-
218 391 26 0 11 
0 0 0 0 0 0 0 0 0 0 
1 0 0
0 0 -8000 0
1 C
3 -26 10 -18
0
0
0
24 *Combine
*TRAN -1.1 1.1
0
1

0 0 
0 0 0 0 0 0 0 0
0
4441 0 0 0
5 SAVE-
218 179 107 0 11 
0 0 0 0 0 0 0 0 0 0 
1 0 0
0 0 -8000 0
1 B
3 -26 10 -18
0
0
0
10 *TRAN 5u 5
0
1

0 0 
0 0 0 0 0 0 0 0
0
3618 0 0 0
5 SAVE-
218 86 34 0 11 
0 0 0 0 0 0 0 0 0 0 
1 0 0
0 0 -8000 0
1 A
3 -26 10 -18
0
0
0
16 *TRAN -999m 999m
0
1

0 0 
0 0 0 0 0 0 0 0
0
6153 0 0 0
11 Multimeter~
205 532 64 0 22 
0 5 10 11 2 0 0 0 0 0 
78 79 32 68 65 84 65 32 0 0 
0 82 0 0
0 0 16448 0
8 1.000Meg
-28 -19 28 -11
4 R0m1
-14 -29 14 -21
0
0
11 %D %1 %4 %V
0
5

0 1 2 3 4 0 
82 0 0 0 0 0 0 0
1 R
5394 0 0 0
2 +V
167 479 21 0 2 
0 6 0 0
0 0 -11424 0
2 5V
8 -3 22 5
2 V1
7 -13 21 -5
0
0
13 %D %1 0 DC %V
0
2

0 1 0 
86 0 0 0 0 0 0 0
1 V
7734 0 0 0
7 Ground~
168 409 138 0 2 
0 2 0 0
0 0 -12192 0
0
0
0
4 GND;
0
0
2

0 1 0 
0 0 0 0 0 0 0 0
0
9914 0 0 0
11 Signal Gen~
195 350 41 0 -15 
0 4 2 2 86 -8 8 0 0 0 
0 0 0 0 0 0 
1.000000 1000000.000000 0.000000 1.100000 0.000000 
0.000000 0.000000 0.000000 0.000000 0.000000 
0.000000 0.000000 0.000000 0.000000 0.000000 
0.000000 0.000000 0.000000 0.000000 0.000000 0
0 0 16960 0
5 -1/1V
-15 -48 20 -40
2 V2
-8 -32 6 -24
0
0
40 %D %1 %2 DC 0 SIN(0 1.1 1Meg 0 0) AC 1 0
0
3

0 1 2 0 
86 0 0 0 0 0 0 0
1 V
3747 0 0 0
10 I->Switch~
94 459 69 0 5 
0 6 5 3 2 0 10 I->Switch~
1 0 576 0
3 CSW
-24 -37 -3 -29
5 IcSw1
-17 12 18 20
0
0
32 V%D %3 %4 DC 0V
%D %1 %2 V%D %M
0
5

0 3 4 1 2 0 
87 0 0 0 0 0 0 0
4 IcSw
3549 0 0 0
11 Multimeter~
205 204 68 0 22 
0 7 12 13 2 0 0 0 0 0 
78 79 32 68 65 84 65 32 0 0 
0 82 0 0
0 0 16448 0
8 1.000Meg
-28 -19 28 -11
4 R0m2
-14 -29 14 -21
0
0
11 %D %1 %4 %V
0
5

0 1 2 3 4 0 
82 0 0 0 0 0 0 0
1 R
7931 0 0 0
7 Ground~
168 97 156 0 2 
0 2 0 0
0 0 -12192 0
0
0
0
4 GND;
0
0
2

0 1 0 
0 0 0 0 0 0 0 0
0
9325 0 0 0
11 Signal Gen~
195 39 39 0 -15 
0 8 2 2 86 -10 10 0 0 0 
0 0 0 0 0 0 
0.000000 1000000.000000 0.000000 1.000000 0.000000 
0.000000 0.000000 0.000000 0.000000 0.000000 
0.000000 0.000000 0.000000 0.000000 0.000000 
0.000000 0.000000 0.000000 0.000000 0.000000 0
0 0 16960 0
5 -1/1V
-15 -48 20 -40
2 V3
-7 -30 7 -22
0
0
31 %D %1 %2 DC 0 SIN(0 1 1Meg 0 0)
0
3

0 1 2 0 
86 0 0 0 0 0 0 0
1 V
8903 0 0 0
2 +V
167 137 17 0 2 
0 9 0 0
0 0 -11424 0
2 5V
6 5 20 13
2 V4
7 -6 21 2
0
0
13 %D %1 0 DC %V
0
2

0 1 0 
86 0 0 0 0 0 0 0
1 V
3834 0 0 0
10 V->Switch~
94 117 69 0 5 
0 9 7 8 2 0 10 V->Switch~
2 0 576 0
4 SW05
-14 -37 14 -29
5 VcIs1
-17 12 18 20
0
0
17 %D %1 %2 %3 %4 %M
0
5

0 3 4 1 2 0 
83 0 0 0 0 0 0 0
4 VcIs
3363 0 0 0
9 Resistor~
94 416 26 0 3 
0 4 3 0 9 Resistor~
3 0 4960 0
2 1k
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
3

0 1 2 0 
82 0 0 0 0 0 0 0
1 R
7668 0 0 0
13
2 3 3 0 0 8320 0 15 9 0 0 3
434 26
439 26
439 42
1 1 4 0 0 12416 0 8 15 0 0 4
381 36
387 36
387 26
398 26
4 0 2 0 0 8320 0 5 0 0 7 3
557 87
557 120
409 120
2 1 5 0 0 8320 0 9 5 0 0 4
479 96
479 106
507 106
507 87
1 1 6 0 0 12416 0 6 9 0 0 4
479 30
479 27
479 27
479 42
4 0 2 0 0 0 0 9 0 0 7 3
439 96
439 107
409 107
2 1 2 0 0 0 0 8 7 0 0 3
381 46
409 46
409 132
1 2 7 0 0 8320 0 10 14 0 0 4
179 91
179 122
137 122
137 96
4 0 2 0 0 0 0 10 0 0 11 3
229 91
229 137
97 137
2 0 2 0 0 0 0 12 0 0 11 3
70 44
70 137
97 137
4 1 2 0 0 0 0 14 11 0 0 2
97 96
97 150
1 3 8 0 0 4224 0 12 14 0 0 3
70 34
97 34
97 42
1 1 9 0 0 4224 0 13 14 0 0 2
137 26
137 42
0
0
17 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2.5e-008 2.5e-008 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
