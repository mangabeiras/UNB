CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 27 100 9
16 74 624 456
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
16 74 624 456
145227798 0
0
0
0
0
0
0
4
7 Ground~
168 266 210 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
8 Battery~
219 163 148 0 2 64
0 7 2
8 Battery~
0 0 320 0
3 10V
12 -5 33 3
2 V1
15 -15 29 -7
0
0
14 %D %1 %2 DC %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 1 0 0
1 V
4441 0 0
0
0
9 Resistor~
219 224 108 0 2 64
0 7 6
9 Resistor~
0 0 352 0
2 1k
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
9 Resistor~
219 319 108 0 4 64
0 6 2 0 -1
9 Resistor~
0 0 352 0
2 1k
-7 -12 7 -4
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
7
0 0 3 0 0 4224 0 0 0 0 0 3
224 116
224 139
241 139
0 0 4 0 0 4224 0 0 0 0 0 3
179 102
179 39
239 39
0 0 5 0 0 4224 0 0 0 0 0 3
210 101
210 63
240 63
2 1 6 0 0 4224 0 3 4 0 0 2
242 108
301 108
1 1 7 0 0 8320 0 2 3 0 0 3
163 135
163 108
206 108
1 0 2 0 0 4096 0 1 0 0 7 2
266 204
266 190
2 2 2 0 0 12416 0 4 2 0 0 5
337 108
359 108
359 190
163 190
163 159
3
-11 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 39
243 128 331 182
247 132 328 174
39 Measure power
dissipation on a
device
-11 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 24
241 52 363 72
245 56 360 70
24 Measure current on a pin
-11 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 25
241 28 368 48
245 32 365 46
25 Measure voltage on a wire
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
