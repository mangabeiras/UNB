CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
0 66 640 259
144179216 0
0
0
0
0
0
0
8
5 SAVE-
218 164 38 0 64 64
0 0 0 0 0 0 0 0 0 0
1 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -1610612472
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
16 *DC -435p 3.49 0
0
0
0
1

0 0
0 0 0 0 1 0 0 0
4 SAVE
8953 0 0
0
0
7 Ground~
168 33 73 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 261 74 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
9 V Source~
197 162 56 0 2 5
0 4 3
0
0 0 16736 0
2 0V
15 -2 29 6
2 V1
15 -12 29 -4
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
6153 0 0
0
0
9 V Source~
197 214 56 0 2 5
0 2 3
0
0 0 16992 0
3 10V
12 -2 33 6
3 VDS
12 -12 33 -4
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
5394 0 0
0
0
9 V Source~
197 70 75 0 2 5
0 2 5
0
0 0 16992 0
3 10V
12 -2 33 6
3 VGS
12 -12 33 -4
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
7734 0 0
0
0
7 Ground~
168 133 123 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
12 P-EMOS 3T:A~
219 127 92 0 3 7
0 4 5 2
12 P-EMOS 3T:A~
0 0 832 0
7 IRF9510
16 8 65 16
3 Q1A
30 -3 51 5
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-220
7

0 2 1 3 2 1 3 -33686019
109 0 552 256 1 1 0 0
1 Q
3747 0 0
0
0
6
2 2 3 0 0 8320 0 4 5 0 0 4
162 77
162 84
214 84
214 77
1 1 4 0 0 4224 0 8 4 0 0 4
133 74
133 28
162 28
162 35
1 1 2 0 0 8320 0 3 5 0 0 4
261 68
261 28
214 28
214 35
1 1 2 0 0 0 0 6 2 0 0 4
70 54
70 47
33 47
33 67
2 2 5 0 0 8320 0 6 8 0 0 3
70 96
70 101
109 101
3 1 2 0 0 0 0 8 7 0 0 2
133 110
133 117
0
0
4 0 0
0
0
3 VDS
0 15 0.1
3 VGS
5 10 1
3 0 1 4
0 8e-007 1e-008 1e-008 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
1520 2259520 100 100 0 0
98 66 608 126
0 259 640 452
608 66
98 66
608 66
608 126
0 0
5.43943e-315 5.2221e-315 5.5705e-315 0 5.43813e-315 5.5705e-315
12409 0
4 3 10
1
162 38
0 4 0 0 1	4 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
