CircuitMaker Text
5.6
Probes: 2
V1_1
Transient Analysis
0 107 102 65280
LLTR1_3
Transient Analysis
1 224 103 65535
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
245 80 925 597
7 5.000 V
7 5.000 V
3 GND
5e+07 10
24 100 0 1 0
20 Package,Description,
64 D:\Program Files\Protel Technology\CircuitMaker 2000 Pro\BOM.DAT
0 7
2 4 0.500000 0.500000
245 339 925 597
9961474 0
0
0
0
0
0
0
5
7 Ground~
168 248 137 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
7422 0 0
2
36626.4 0
0
7 Ground~
168 111 136 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3557 0 0
2
36626.4 1
0
11 Signal Gen~
195 64 106 0 24 64
0 4 2 1 86 -9 9 0 0 0
0 0 0 0 0 0 0 1268291200 0 1084227584
0 822702175 822702175 850119799 861323157
20
0 2e+07 0 5 0 2e-09 2e-09 2e-08 5e-08 0
0 0 0 0 0 0 0 0 0 0
0
0 0 16976 0
5 -1/1V
-15 -48 20 -40
2 V1
-6 -35 8 -27
0
0
40 %D %1 %2 DC 0 PULSE(0 5 0 2n 2n 20n 50n)
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
3459 0 0
2
36626.4 2
0
13 LossLessLine~
219 173 107 0 4 64
0 4 2 3 2
13 LossLessLine~
0 0 848 0
13 ZO=50 TD=20NS
-46 -20 45 -12
5 LLTR1
-18 -30 17 -22
0
0
17 %D %1 %2 %3 %4 %L
0
0
0
9

0 1 2 3 4 1 2 3 4 -33686019
84 0 0 0 1 0 0 0
4 LLTR
3684 0 0
2
36626.4 3
0
9 Resistor~
219 245 103 0 4 64
0 3 2 0 -1
9 Resistor~
0 0 4976 0
2 1k
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
9470 0 0
2
36626.4 4
0
6
1 0 2 0 0 4096 0 2 0 0 5 2
111 130
111 111
1 0 2 0 0 4096 0 1 0 0 4 2
248 131
248 111
1 3 3 0 0 4224 0 5 4 0 0 2
227 103
221 103
4 2 2 0 0 4224 0 4 5 0 0 4
221 111
272 111
272 103
263 103
2 2 2 0 0 0 0 3 4 0 0 2
95 111
125 111
1 1 4 0 0 4224 0 4 3 0 0 4
125 103
100 103
100 101
95 101
0
0
16 0 0
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 1e-07 1e-09 1e-09
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3076 8550464 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
4.29695e-315 0 5.4086e-315 1.60186e-314 4.29695e-315 4.29695e-315
16 0
4 3e-08 5
1
224 103
0 3 0 0 1	0 3 0 0
0 0 100 100 0 0
98 66 294 126
0 0 0 0
294 66
98 66
294 66
294 126
0 0
6.22475e-315 5.26354e-315 5.40943e-315 5.40943e-315 6.22475e-315 6.22475e-315
12403 0
0 3e+06 5e+06
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
5.7175e-315 5.26354e-315 5.31245e-315 0 5.71746e-315 5.71746e-315
16 0
0 500 1000
0
0 0 100 100 0 0
98 66 296 126
0 0 0 0
296 66
98 66
296 66
296 126
0 0
6.08861e-315 5.26354e-315 1.38842e-314 1.38842e-314 6.08861e-315 6.08861e-315
12403 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
