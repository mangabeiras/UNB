CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
50 0 30 100 9
0 66 320 452
7 5.000 V
7 5.000 V
3 GND
2500 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 320 452
9961474 0
0
0
0
0
0
0
12
5 SAVE-
218 310 92 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
30 *Combine
*TRAN -80.00m 80.80m
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 102 117 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
26 *Combine
*TRAN -80m 80.8m
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
2 +V
167 217 27 0 1 64
0 8
0
0 0 54112 0
3 25V
-10 -13 11 -5
2 V1
-6 -24 8 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
7 Ground~
168 164 254 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
11 Signal Gen~
195 53 122 0 19 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1017370378
20
1 1000 0 0.02 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
8 40MV P-P
-28 23 28 31
2 V2
-8 -30 6 -22
0
0
38 %D %1 %2 DC 0 SIN(0 20m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
7 N-JFET~
219 209 117 0 3 64
0 4 5 7
7 N-JFET~
0 0 832 0
6 2N4393
13 -3 55 5
2 Q1
27 -13 41 -5
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 2 3 1 2 3 1 -33686019
74 0 0 0 1 1 0 0
1 Q
7734 0 0
0
0
10 Polar Cap~
219 139 117 0 2 64
0 6 5
10 Polar Cap~
0 0 832 0
3 1uF
-12 -18 9 -10
2 C1
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
10 Polar Cap~
219 289 93 0 2 64
0 4 3
10 Polar Cap~
0 0 832 0
3 1uF
-12 -18 9 -10
2 C2
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
9 Resistor~
219 324 171 0 3 64
0 2 3 -1
9 Resistor~
0 0 4960 90
4 1MEG
5 1 33 9
2 R1
9 -12 23 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 217 181 0 3 64
0 2 7 -1
9 Resistor~
0 0 4960 90
3 500
8 1 29 9
2 R2
9 -12 23 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 217 65 0 4 64
0 4 8 0 1
9 Resistor~
0 0 4960 90
4 2.5K
7 0 35 8
2 R3
9 -12 23 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 164 182 0 3 64
0 2 5 -1
9 Resistor~
0 0 4960 90
4 1MEG
4 -1 32 7
2 R4
11 -13 25 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
12
1 0 2 0 0 8192 0 9 0 0 4 3
324 189
324 233
217 233
2 2 3 0 0 8320 0 8 9 0 0 3
295 93
324 93
324 153
1 0 4 0 0 4224 0 8 0 0 12 2
278 93
217 93
1 2 2 0 0 8320 0 10 5 0 0 5
217 199
217 233
89 233
89 127
84 127
1 0 2 0 0 0 0 4 0 0 6 2
164 248
164 232
1 0 2 0 0 0 0 12 0 0 4 2
164 200
164 233
2 0 5 0 0 4096 0 12 0 0 8 2
164 164
164 117
2 2 5 0 0 4224 0 7 6 0 0 2
145 117
196 117
1 1 6 0 0 4224 0 5 7 0 0 2
84 117
128 117
3 2 7 0 0 4224 0 6 10 0 0 2
217 135
217 163
1 2 8 0 0 4224 0 3 11 0 0 2
217 36
217 47
1 1 4 0 0 0 0 6 11 0 0 2
217 99
217 83
0
0
24 0 0
0
0
0
0 0 0
0
0 0 0
100 0 1 1e+007
0 0.002 1e-005 1e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1432 8550464 100 100 0 0
77 66 287 126
320 66 640 259
286 66
77 66
287 66
287 126
0 0
0 0 0 0 0 0
16 0
4 0.0005 10
2
103 117
0 6 0 0 1	0 9 0 0
324 119
0 3 0 0 2	0 2 0 0
1844 4421696 100 100 0 0
98 66 294 126
320 259 640 452
294 66
98 66
294 66
294 66
0 0
0 0 0 0 0 0
12403 0
4 3e+006 5e+006
1
324 113
0 3 0 0 2	0 2 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
