CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 300 100 3
0 66 645 428
7 5.000 V
7 5.000 V
3 GND
0 66 645 428
9961490 0
0
0
0
0
0
0
53
5 SAVE-
218 683 229 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
20 *Combine
*TRAN -3 3
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 58 129 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
20 *Combine
*TRAN -3 3
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
6 Input~
177 122 419 0 17 64
0 3 0 0 0 0 0 0 0 0
78 70 66 32 32 32 32 32
0
0 0 53344 0
0
0
0
0
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
7 Output~
178 711 186 0 17 64
0 3 0 0 0 0 0 0 0 0
78 70 66 32 32 32 32 32
0
0 0 53344 0
0
0
0
0
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
7 Ground~
168 67 167 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
11 Signal Gen~
195 32 134 0 19 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 0 1148846080 0 1069547520
20
0 1000 0 1.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 16704 0
9 -1.5/1.5V
-31 -28 32 -20
2 V1
-7 -38 7 -30
0
0
31 %D %1 %2 DC 0 SIN(0 1.5 1k 0 0)
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
2 +V
167 578 370 0 1 64
0 4
0
0 0 53600 -19276
5 +420V
7 -10 42 -2
2 V2
17 -20 31 -12
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
2 +V
167 562 394 0 1 64
0 14
0
0 0 53600 -19276
5 +300V
8 -10 43 -2
2 V3
18 -20 32 -12
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
7 Ground~
168 184 281 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
7 Ground~
168 319 244 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
7 Ground~
168 682 295 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
7 Ground~
168 537 262 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
7 Ground~
168 238 428 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
7 Ground~
168 117 389 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
7 Ground~
168 43 247 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
7668 0 0
0
0
2 +V
167 417 227 0 1 64
0 12
0
0 0 53600 90
6 -22.5V
-24 -16 18 -8
2 V4
-4 5 10 13
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
8 Tetrode~
219 128 234 0 4 64
0 28 27 29 7
8 Tetrode~
0 0 320 0
5 7199P
-1 24 34 32
2 Q1
9 14 23 22
0
0
17 %D %1 %2 %3 %4 %S
0
0
0
9

0 1 2 3 4 1 2 3 4 -33686019
88 0 0 0 1 0 0 0
1 Q
3874 0 0
0
0
8 Tetrode~
219 509 290 0 4 64
0 15 14 18 13
8 Tetrode~
0 0 320 -18764
5 6L6GC
10 17 45 25
2 Q2
20 7 34 15
0
0
17 %D %1 %2 %3 %4 %S
0
0
0
9

0 1 2 3 4 1 2 3 4 -33686019
88 0 0 0 1 0 0 0
1 Q
6671 0 0
0
0
8 Tetrode~
219 509 171 0 4 64
0 22 14 23 13
8 Tetrode~
0 0 320 0
5 6L6GC
9 19 44 27
2 Q3
19 9 33 17
0
0
17 %D %1 %2 %3 %4 %S
0
0
0
9

0 1 2 3 4 1 2 3 4 -33686019
88 0 0 0 1 0 0 0
1 Q
3789 0 0
0
0
7 Triode~
219 249 180 0 3 64
0 26 28 9
7 Triode~
0 0 320 0
5 7199T
-3 26 32 34
2 Q4
7 16 21 24
0
0
14 %D %1 %2 %3 %S
0
0
0
7

0 1 2 3 1 2 3 -33686019
88 0 0 0 1 0 0 0
1 Q
4871 0 0
0
0
7 Triode~
219 352 106 0 3 64
0 25 21 20
7 Triode~
0 0 320 0
4 6SN7
1 22 29 30
2 Q5
8 12 22 20
0
0
14 %D %1 %2 %3 %S
0
0
0
7

0 1 2 3 1 2 3 -33686019
88 0 0 0 1 0 0 0
1 Q
3750 0 0
0
0
7 Triode~
219 352 363 0 3 64
0 16 8 19
7 Triode~
0 0 320 -18764
4 6SN7
0 -38 28 -30
2 Q6
7 -48 21 -40
0
0
14 %D %1 %2 %3 %S
0
0
0
7

0 1 2 3 1 2 3 -33686019
88 0 0 0 1 0 0 0
1 Q
8778 0 0
0
0
10 Polar Cap~
219 185 254 0 2 64
0 27 2
10 Polar Cap~
0 0 320 26894
6 0.22uF
5 10 47 18
2 C1
19 0 33 8
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
538 0 0
0
0
10 Capacitor~
219 282 106 0 2 64
0 26 21
10 Polar Cap~
0 0 320 7168
5 0.2uF
-15 -19 20 -11
2 C2
-5 -29 9 -21
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
6843 0 0
0
0
10 Polar Cap~
219 421 62 0 2 64
0 25 24
10 Polar Cap~
0 0 320 7168
5 0.5uF
-19 -18 16 -10
2 C3
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3136 0 0
0
0
10 Polar Cap~
219 422 409 0 2 64
0 16 17
10 Polar Cap~
0 0 320 7168
5 0.5uF
-18 14 17 22
2 C4
-8 8 6 16
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
5950 0 0
0
0
10 Polar Cap~
219 274 357 0 2 64
0 9 8
10 Polar Cap~
0 0 320 7168
5 0.2uF
-12 12 23 20
2 C5
-2 2 12 10
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
5670 0 0
0
0
14 CTTransformer~
219 623 243 0 5 64
0 3 2 22 4 15
14 CTTransformer~
0 0 64 512
0
2 T1
-7 -40 7 -32
0
0
104 LA%D %1 %2 0.01
LB%D %3 %4 2.2
LC%D %4 %5 2.2
%DA LA%D LB%D .99
%DB LA%D LC%D .99
%DC LB%D LC%D .99
0
0
0
11

0 1 2 3 4 5 1 2 3 4
5 -33686019
75 0 0 0 1 0 0 0
1 T
6828 0 0
0
0
9 Resistor~
219 88 208 0 2 64
0 29 5
9 Resistor~
0 0 352 90
3 10k
6 -5 27 3
2 R1
9 -15 23 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 43 207 0 3 64
0 2 5 -1
9 Resistor~
0 0 352 90
4 100k
4 -5 32 3
2 R2
11 -15 25 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 128 100 0 4 64
0 28 14 0 1
9 Resistor~
0 0 352 90
4 220k
-36 -8 -8 0
2 R3
-29 -18 -15 -10
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 184 101 0 4 64
0 27 14 0 1
9 Resistor~
0 0 352 90
4 820k
9 -5 37 3
2 R4
16 -15 30 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
9 Resistor~
219 249 76 0 4 64
0 26 14 0 1
9 Resistor~
0 0 352 90
3 15k
-27 -3 -6 5
2 R5
-24 -13 -10 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3635 0 0
0
0
9 Resistor~
219 387 94 0 3 64
0 4 25 1
9 Resistor~
0 0 352 90
3 47k
6 -2 27 6
2 R6
6 -11 20 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3973 0 0
0
0
9 Resistor~
219 438 89 0 3 64
0 12 24 1
9 Resistor~
0 0 352 90
4 100k
4 -4 32 4
2 R7
6 -14 20 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3851 0 0
0
0
9 Resistor~
219 473 145 0 2 64
0 23 24
9 Resistor~
0 0 352 90
4 3.9k
4 -5 32 3
2 R8
6 -14 20 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8383 0 0
0
0
9 Resistor~
219 682 243 0 3 64
0 2 3 -1
9 Resistor~
0 0 352 90
1 8
9 -2 16 6
2 R9
6 -12 20 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
9 Resistor~
219 117 292 0 2 64
0 6 7
9 Resistor~
0 0 352 90
3 820
7 -2 28 6
3 R10
7 -12 28 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 117 351 0 3 64
0 2 6 -1
9 Resistor~
0 0 352 90
2 22
5 -2 19 6
3 R11
2 -12 23 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3334 0 0
0
0
9 Resistor~
219 169 353 0 2 64
0 3 6
9 Resistor~
0 0 352 90
3 390
6 -3 27 5
3 R12
6 -13 27 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3559 0 0
0
0
9 Resistor~
219 238 392 0 3 64
0 2 9 -1
9 Resistor~
0 0 352 90
3 15k
8 -2 29 6
3 R13
8 -12 29 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
984 0 0
0
0
9 Resistor~
219 304 320 0 2 64
0 8 10
9 Resistor~
0 0 352 90
4 1Meg
-33 -4 -5 4
3 R14
3 -14 24 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7557 0 0
0
0
9 Resistor~
219 341 301 0 2 64
0 19 10
9 Resistor~
0 0 352 90
2 1k
7 -3 21 5
3 R15
4 -13 25 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3146 0 0
0
0
9 Resistor~
219 341 250 0 4 64
0 10 2 0 -1
9 Resistor~
0 0 352 90
4 3.8k
5 -4 33 4
3 R16
3 -14 24 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
5687 0 0
0
0
9 Resistor~
219 341 156 0 2 64
0 11 20
9 Resistor~
0 0 352 90
2 1k
6 -3 20 5
3 R17
3 -13 24 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7939 0 0
0
0
9 Resistor~
219 341 200 0 3 64
0 2 11 -1
9 Resistor~
0 0 352 90
4 3.8k
6 -4 34 4
3 R18
3 -16 24 -8
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3308 0 0
0
0
9 Resistor~
219 307 136 0 2 64
0 11 21
9 Resistor~
0 0 352 90
4 1Meg
-32 -3 -4 5
3 R19
4 -12 25 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3408 0 0
0
0
9 Resistor~
219 408 310 0 2 64
0 15 10
9 Resistor~
0 0 352 90
3 75k
5 -6 26 2
3 R20
2 -12 23 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
9773 0 0
0
0
9 Resistor~
219 387 370 0 4 64
0 16 4 0 1
9 Resistor~
0 0 352 90
3 47k
7 -5 28 3
3 R21
3 -14 24 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
691 0 0
0
0
9 Resistor~
219 438 370 0 4 64
0 17 12 0 1
9 Resistor~
0 0 352 90
4 100k
5 -2 33 6
3 R22
4 -15 25 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7834 0 0
0
0
9 Resistor~
219 474 311 0 2 64
0 17 18
9 Resistor~
0 0 352 90
4 3.9k
4 -3 32 5
3 R23
3 -15 24 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3588 0 0
0
0
9 Resistor~
219 408 148 0 2 64
0 11 22
9 Resistor~
0 0 352 90
3 75k
5 -4 26 4
3 R24
2 -14 23 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4528 0 0
0
0
9 Resistor~
219 537 226 0 3 64
0 2 13 -1
9 Resistor~
0 0 352 90
2 10
6 -5 20 3
3 R25
3 -15 24 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3303 0 0
0
0
65
0 0 4 0 0 4096 0 0 0 4 2 2
578 251
387 251
1 2 4 0 0 4224 0 34 49 0 0 2
387 112
387 352
2 0 2 0 0 12416 0 28 0 0 30 4
642 251
650 251
650 272
682 272
4 1 4 0 0 0 0 28 7 0 0 3
604 243
578 243
578 355
1 0 3 0 0 8192 0 4 0 0 31 3
671 186
663 186
663 221
1 1 3 0 0 8320 0 3 40 0 0 3
156 419
169 419
169 371
2 1 2 0 0 0 0 6 5 0 0 3
63 139
67 139
67 161
1 0 5 0 0 8320 0 6 0 0 9 3
63 129
81 129
81 182
2 2 5 0 0 0 0 30 29 0 0 4
43 189
43 182
88 182
88 190
2 0 6 0 0 8320 0 40 0 0 12 3
169 335
169 316
117 316
1 1 2 0 0 0 0 39 14 0 0 2
117 369
117 383
1 2 6 0 0 0 0 38 39 0 0 2
117 310
117 333
2 4 7 0 0 4224 0 38 17 0 0 2
117 274
117 257
1 0 8 0 0 4096 0 42 0 0 15 2
304 338
304 357
2 2 8 0 0 4224 0 27 22 0 0 2
280 357
326 357
1 0 9 0 0 4096 0 27 0 0 18 2
263 357
238 357
1 1 2 0 0 0 0 41 13 0 0 2
238 410
238 422
3 2 9 0 0 4224 0 20 41 0 0 2
238 203
238 374
2 0 10 0 0 8192 0 42 0 0 22 3
304 302
304 277
341 277
1 0 11 0 0 8192 0 47 0 0 23 3
307 154
307 177
341 177
0 1 2 0 0 0 0 0 10 41 0 3
341 224
319 224
319 238
2 0 10 0 0 8320 0 48 0 0 40 3
408 292
408 277
341 277
1 0 11 0 0 8320 0 52 0 0 42 3
408 166
408 177
341 177
1 0 12 0 0 4096 0 16 0 0 45 2
428 225
438 225
2 0 13 0 0 8192 0 53 0 0 28 3
537 208
537 201
498 201
1 1 2 0 0 0 0 12 53 0 0 2
537 256
537 244
2 0 14 0 0 4096 0 18 0 0 29 2
535 287
562 287
4 4 13 0 0 4224 0 19 18 0 0 2
498 194
498 261
2 1 14 0 0 8192 0 19 8 0 0 3
535 168
562 168
562 379
1 1 2 0 0 0 0 37 11 0 0 2
682 261
682 289
2 1 3 0 0 0 0 37 28 0 0 5
682 225
682 221
650 221
650 235
642 235
1 0 15 0 0 4096 0 18 0 0 33 2
509 310
509 333
1 5 15 0 0 8320 0 48 28 0 0 5
408 328
408 333
593 333
593 259
604 259
1 0 16 0 0 4096 0 49 0 0 38 2
387 388
387 409
1 0 17 0 0 4096 0 50 0 0 36 2
438 388
438 409
1 2 17 0 0 4224 0 51 26 0 0 3
474 329
474 409
428 409
3 2 18 0 0 8320 0 18 51 0 0 3
483 281
474 281
474 293
1 1 16 0 0 8320 0 22 26 0 0 3
352 383
352 409
411 409
1 3 19 0 0 4224 0 43 22 0 0 2
341 319
341 334
1 2 10 0 0 0 0 44 43 0 0 2
341 268
341 283
1 2 2 0 0 0 0 46 44 0 0 2
341 218
341 232
1 2 11 0 0 0 0 45 46 0 0 2
341 174
341 182
3 2 20 0 0 4224 0 21 45 0 0 2
341 129
341 138
2 0 21 0 0 4096 0 47 0 0 54 2
307 118
307 106
1 2 12 0 0 4224 0 35 50 0 0 2
438 107
438 352
1 0 22 0 0 4096 0 19 0 0 47 2
509 145
509 118
2 3 22 0 0 8320 0 52 28 0 0 5
408 130
408 118
593 118
593 227
604 227
1 3 23 0 0 4224 0 36 19 0 0 3
473 163
473 174
483 174
2 0 24 0 0 4096 0 35 0 0 50 2
438 71
438 62
2 2 24 0 0 4224 0 36 25 0 0 3
473 127
473 62
427 62
2 0 25 0 0 4096 0 34 0 0 52 2
387 76
387 62
1 1 25 0 0 4224 0 25 21 0 0 3
410 62
352 62
352 80
1 0 26 0 0 4096 0 24 0 0 56 2
271 106
249 106
2 2 21 0 0 4224 0 24 21 0 0 2
288 106
326 106
2 0 14 0 0 0 0 33 0 0 62 2
249 58
249 37
1 1 26 0 0 4224 0 20 33 0 0 2
249 154
249 94
2 0 27 0 0 4096 0 17 0 0 60 2
154 231
184 231
2 0 14 0 0 0 0 32 0 0 62 2
184 83
184 37
2 1 2 0 0 0 0 23 9 0 0 2
184 261
184 275
1 1 27 0 0 4224 0 32 23 0 0 2
184 119
184 244
2 0 28 0 0 4224 0 20 0 0 63 2
223 180
128 180
2 0 14 0 0 8320 0 31 0 0 29 4
128 82
128 37
562 37
562 168
1 1 28 0 0 0 0 17 31 0 0 2
128 208
128 118
1 3 29 0 0 8320 0 29 17 0 0 3
88 226
88 237
102 237
1 1 2 0 0 0 0 30 15 0 0 2
43 225
43 241
1
-16 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 27
256 4 536 33
260 8 530 27
27 Vacuum-tube Power Amplifier
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.005 2.5e-005 2.5e-005 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
1544 1210432 100 100 0 0
0 0 0 0
0 60 140 130
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
4 1 200
0
1548 8550464 100 100 0 0
77 66 977 276
0 401 1024 742
977 66
77 66
977 66
977 276
0 0
4.94359e-315 0 5.44981e-315 1.60615e-314 4.94359e-315 5.49213e-315
16 0
4 0.001 300
1
669 221
0 3 0 0 2	0 31 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
