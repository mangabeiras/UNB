CircuitMaker Text
5.6
Probes: 17
U6A_3
AC Analysis
2 246 254 16776960
U6A_3
DC Sweep
2 246 254 16776960
U6A_3
Operating Point
2 246 254 16776960
U6A_3
Fourier Analysis
2 246 254 16776960
U1E_11
AC Analysis
0 302 186 65280
U1E_11
DC Sweep
0 302 186 65280
U1E_11
Operating Point
0 302 186 65280
U1E_11
Fourier Analysis
0 302 186 65280
U5A_1
AC Analysis
1 200 165 65535
U5A_1
DC Sweep
1 200 165 65535
U5A_1
Operating Point
1 200 165 65535
U5A_1
Fourier Analysis
1 200 165 65535
Clk
Transient Analysis
0 201 159 65280
Q0
Transient Analysis
1 514 186 65535
Q1
Transient Analysis
2 514 230 16776960
Q2
Transient Analysis
3 514 274 16711935
Q3
Transient Analysis
4 536 309 11184640
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 80 3 80 10
231 152 911 669
7 5.000 V
7 5.000 V
3 GND
100000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
2 4 0.500000 0.500000
231 411 911 669
11010054 0
0
0
0
0
0
0
33
13 Logic Switch~
5 154 271 0 1 11
0 8
0
0 0 4464 0
2 0V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9496 0 0
2
5.8901e-315 0
0
13 Logic Switch~
5 156 298 0 1 11
0 9
0
0 0 4464 0
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5392 0 0
2
5.8901e-315 5.26354e-315
0
9 Inverter~
13 580 324 0 2 21
0 7 16
0
0 0 112 0
4 4069
-14 -19 14 -11
3 U4B
-11 -29 10 -21
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 2 4 0
1 U
3710 0 0
2
5.8901e-315 5.32571e-315
0
9 Inverter~
13 577 274 0 2 21
0 6 15
0
0 0 112 0
4 4069
-14 -19 14 -11
3 U4A
-11 -29 10 -21
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 1 4 0
1 U
6540 0 0
2
5.8901e-315 5.34643e-315
0
9 Inverter~
13 576 230 0 2 21
0 5 14
0
0 0 112 0
4 4069
-14 -19 14 -11
3 U1F
-11 -29 10 -21
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 6 1 0
1 U
9337 0 0
2
5.8901e-315 5.3568e-315
0
9 Inverter~
13 576 186 0 2 21
0 4 13
0
0 0 112 0
4 4069
-14 -19 14 -11
3 U1E
-11 -29 10 -21
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 5 1 0
1 U
5573 0 0
2
5.8901e-315 5.36716e-315
0
10 2-In NAND~
219 213 285 0 3 21
0 8 9 12
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U6A
-4 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 6 0
1 U
6668 0 0
2
5.8901e-315 5.37752e-315
0
6 74112~
219 498 160 0 7 31
0 11 11 6 11 12 25 7
0
0 0 4208 0
7 74LS112
-3 -60 46 -52
3 U3A
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 1 3 0
1 U
4641 0 0
2
5.8901e-315 5.38788e-315
0
6 74112~
219 414 160 0 7 31
0 11 11 5 11 12 26 6
0
0 0 4208 0
7 74LS112
-3 -60 46 -52
3 U2A
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 1 2 0
1 U
6837 0 0
2
5.8901e-315 5.39306e-315
0
6 74112~
219 327 159 0 7 31
0 11 11 4 11 12 27 5
0
0 0 4208 0
7 74LS112
-3 -60 46 -52
3 U5B
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 2 5 0
1 U
3462 0 0
2
5.8901e-315 5.39824e-315
0
6 74112~
219 245 158 0 7 31
0 11 11 3 11 12 28 4
0
0 0 4208 0
7 74LS112
-3 -60 46 -52
3 U5A
11 -70 32 -62
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 -33686019
65 0 0 512 2 1 5 0
1 U
3526 0 0
2
5.8901e-315 5.40342e-315
0
2 +V
167 698 66 0 1 3
0 10
0
0 0 53616 0
4 +15V
-14 -22 14 -14
2 V3
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3159 0 0
2
5.8901e-315 5.41896e-315
0
7 Ground~
168 765 363 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6490 0 0
2
5.8901e-315 5.42414e-315
0
7 Ground~
168 721 308 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7652 0 0
2
5.8901e-315 5.42933e-315
0
7 Ground~
168 675 261 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
954 0 0
2
5.8901e-315 5.43192e-315
0
7 Ground~
168 627 215 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6174 0 0
2
5.8901e-315 5.43451e-315
0
2 +V
167 340 64 0 1 3
0 11
0
0 0 53616 0
3 +5V
-10 -15 11 -7
2 V4
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6578 0 0
2
5.8901e-315 5.4371e-315
0
12 NPN Trans:C~
219 622 186 0 3 7
0 20 13 2
12 NPN Trans:C~
0 0 336 0
3 NPN
17 -5 38 3
2 Q1
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
962 0 0
2
5.8901e-315 5.43969e-315
0
12 NPN Trans:C~
219 670 230 0 3 7
0 19 14 2
12 NPN Trans:C~
0 0 336 0
3 NPN
17 -5 38 3
2 Q2
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
4850 0 0
2
5.8901e-315 5.44228e-315
0
12 NPN Trans:C~
219 716 274 0 3 7
0 18 15 2
12 NPN Trans:C~
0 0 336 0
3 NPN
17 -5 38 3
2 Q3
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
3841 0 0
2
5.8901e-315 5.44487e-315
0
12 NPN Trans:C~
219 760 324 0 3 7
0 17 16 2
12 NPN Trans:C~
0 0 336 0
3 NPN
17 -5 38 3
2 Q4
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 1 0 0
1 Q
8581 0 0
2
5.8901e-315 5.44746e-315
0
4 .IC~
207 24 169 0 1 3
0 23
0
0 0 53584 0
2 0V
-7 -15 7 -7
4 CMD1
-14 -25 14 -17
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
3 CMD
9945 0 0
2
5.8901e-315 5.45005e-315
0
2 +V
167 103 78 0 1 3
0 21
0
0 0 53616 0
3 +5V
-11 -22 10 -14
2 V5
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5593 0 0
2
5.8901e-315 5.45264e-315
0
10 555 Timer~
219 141 143 0 8 17
0 2 23 3 21 22 23 24 21
10 555 Timer~
0 0 6480 0
3 555
-10 -23 11 -15
2 U7
-7 -33 7 -25
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 -33686019
88 0 0 0 1 1 0 0
1 U
7654 0 0
2
5.8901e-315 5.45523e-315
0
10 Polar Cap~
219 52 218 0 2 5
0 23 2
10 Polar Cap~
0 0 848 26894
5 .01uF
-48 2 -13 10
2 C1
-33 -8 -19 0
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
6858 0 0
2
5.8901e-315 5.45782e-315
0
10 Polar Cap~
219 176 213 0 2 5
0 22 2
10 Polar Cap~
0 0 848 26894
5 .01uF
10 4 45 12
2 C2
21 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
3228 0 0
2
5.8901e-315 5.46041e-315
0
7 Ground~
168 90 252 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4179 0 0
2
5.8901e-315 5.463e-315
0
9 Resistor~
219 628 134 0 4 5
0 20 10 0 1
9 Resistor~
0 0 368 90
2 1k
8 -5 22 3
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
9618 0 0
2
5.8901e-315 5.46559e-315
0
9 Resistor~
219 675 137 0 4 5
0 19 10 0 1
9 Resistor~
0 0 368 90
2 1k
8 -5 22 3
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
8659 0 0
2
5.8901e-315 5.46818e-315
0
9 Resistor~
219 721 137 0 4 5
0 18 10 0 1
9 Resistor~
0 0 368 90
2 1k
8 -5 22 3
2 R3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
6117 0 0
2
5.8901e-315 5.47077e-315
0
9 Resistor~
219 765 140 0 4 5
0 17 10 0 1
9 Resistor~
0 0 368 90
2 1k
8 -5 22 3
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
6779 0 0
2
5.8901e-315 5.47207e-315
0
9 Resistor~
219 51 173 0 2 5
0 23 24
9 Resistor~
0 0 4976 90
3 500
4 0 25 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3927 0 0
2
5.8901e-315 5.47336e-315
0
9 Resistor~
219 51 116 0 4 5
0 24 21 0 1
9 Resistor~
0 0 4976 90
3 100
7 0 28 8
2 R6
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
5610 0 0
2
5.8901e-315 5.47466e-315
0
55
0 1 2 0 0 4096 0 0 27 46 0 4
90 235
90 248
90 248
90 246
3 3 3 0 0 12416 0 24 11 0 0 6
109 152
98 152
98 179
200 179
200 131
215 131
1 1 8 0 0 4224 0 1 7 0 0 4
166 271
179 271
179 276
189 276
1 2 9 0 0 12416 0 2 7 0 0 4
168 298
178 298
178 294
189 294
3 0 4 0 0 4096 0 10 0 0 6 2
297 132
283 132
7 1 4 0 0 12416 0 11 6 0 0 4
269 122
283 122
283 186
561 186
1 0 10 0 0 4096 0 12 0 0 36 2
698 75
698 99
1 0 11 0 0 4096 0 10 0 0 21 2
327 96
327 84
7 1 7 0 0 8336 0 8 3 0 0 4
522 124
535 124
535 324
565 324
0 1 6 0 0 4224 0 0 4 22 0 3
451 133
451 274
562 274
1 0 11 0 0 8192 0 8 0 0 21 3
498 97
498 84
459 84
1 0 11 0 0 0 0 9 0 0 21 2
414 97
414 84
1 0 11 0 0 0 0 11 0 0 21 2
245 95
245 84
1 0 11 0 0 0 0 17 0 0 21 2
340 73
340 84
2 0 11 0 0 0 0 8 0 0 21 2
474 124
459 124
2 0 11 0 0 0 0 9 0 0 17 2
390 124
378 124
4 0 11 0 0 8192 0 9 0 0 21 3
390 142
378 142
378 84
2 0 11 0 0 0 0 10 0 0 19 2
303 123
293 123
4 0 11 0 0 0 0 10 0 0 21 3
303 141
293 141
293 84
2 0 11 0 0 0 0 11 0 0 21 2
221 122
210 122
4 4 11 0 0 12416 0 11 8 0 0 6
221 140
210 140
210 84
459 84
459 142
474 142
7 3 6 0 0 0 0 9 8 0 0 4
438 124
451 124
451 133
468 133
5 0 12 0 0 4096 0 9 0 0 43 2
414 172
414 206
5 0 12 0 0 4096 0 10 0 0 43 2
327 171
327 206
2 2 13 0 0 4224 0 18 6 0 0 2
604 186
597 186
2 2 14 0 0 4224 0 5 19 0 0 2
597 230
652 230
2 2 15 0 0 4224 0 20 4 0 0 2
698 274
598 274
2 2 16 0 0 4224 0 3 21 0 0 2
601 324
742 324
1 0 5 0 0 4224 0 5 0 0 41 3
561 230
368 230
368 133
3 1 2 0 0 4096 0 21 13 0 0 2
765 342
765 357
3 1 2 0 0 0 0 20 14 0 0 2
721 292
721 302
3 1 2 0 0 0 0 19 15 0 0 2
675 248
675 255
3 1 2 0 0 0 0 18 16 0 0 2
627 204
627 209
2 0 10 0 0 0 0 30 0 0 36 2
721 119
721 99
2 0 10 0 0 0 0 29 0 0 36 2
675 119
675 99
2 2 10 0 0 8320 0 28 31 0 0 4
628 116
628 99
765 99
765 122
1 1 17 0 0 4224 0 31 21 0 0 2
765 158
765 306
1 1 18 0 0 4224 0 30 20 0 0 2
721 155
721 256
1 1 19 0 0 4224 0 29 19 0 0 2
675 155
675 212
1 1 20 0 0 4224 0 28 18 0 0 4
628 152
628 160
627 160
627 168
7 3 5 0 0 0 0 10 9 0 0 4
351 123
368 123
368 133
384 133
5 0 12 0 0 4096 0 11 0 0 43 2
245 170
245 206
3 5 12 0 0 12416 0 7 8 0 0 5
240 285
245 285
245 206
498 206
498 172
8 1 21 0 0 8192 0 24 23 0 0 3
173 134
173 87
103 87
1 0 2 0 0 8192 0 24 0 0 46 3
109 134
76 134
76 235
2 2 2 0 0 8320 0 26 25 0 0 4
175 220
175 235
51 235
51 225
5 1 22 0 0 8320 0 24 26 0 0 3
173 161
175 161
175 203
1 0 23 0 0 8192 0 22 0 0 49 3
24 181
24 192
51 192
0 0 23 0 0 4096 0 0 0 52 55 2
51 192
91 192
2 1 21 0 0 0 0 33 23 0 0 3
51 98
51 87
103 87
7 0 24 0 0 12416 0 24 0 0 53 6
173 143
188 143
188 112
86 112
86 143
51 143
1 1 23 0 0 0 0 32 25 0 0 2
51 191
51 208
1 2 24 0 0 0 0 33 32 0 0 2
51 134
51 155
4 1 21 0 0 8320 0 24 23 0 0 3
109 161
103 161
103 87
2 6 23 0 0 12416 0 24 24 0 0 6
109 143
91 143
91 192
186 192
186 152
173 152
6
-20 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 40
171 22 660 57
175 26 655 53
40 Mixed-mode Binary Ripple Counter Circuit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 3
200 163 226 178
200 163 226 178
3 Clk
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
546 171 564 186
546 171 564 186
2 Q0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
545 215 563 230
545 215 563 230
2 Q1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
547 259 565 274
547 259 565 274
2 Q2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
548 309 566 324
548 309 566 324
2 Q3
33 .OPTIONS ITL4=100.0 TRTOL=3.000

16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.0001 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2492 8526400 100 100 0 0
98 66 608 126
0 259 640 452
608 66
98 66
608 66
608 126
0 0
0 0 0 0 0 0
12409 0
4 1e-05 10
1
619 161
0 20 0 0 1	0 40 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
