CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 18 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 800 319
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 800 319
10027026 0
0
6 Title:
5 Name:
0
0
0
5
4 DAC8
219 171 83 0 11 23
0 12 11 10 9 8 7 6 5 2
4 3
4 DAC8
0 0 13040 0
4 DAC8
-14 -55 14 -47
2 U1
-7 -55 7 -47
0
16 DVCC=14;DGND=13;
108 %D [%14bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %11o] %M
0
12 type:digital
5 DIP14
23

0 1 2 3 4 5 6 7 8 9
10 11 1 2 3 4 5 6 7 8
9 10 11 0
65 0 0 0 1 0 0 0
1 U
8953 0 0
0
0
9 Data Seq~
170 51 83 0 17 18
0 12 11 10 9 8 7 6 5 13
14 1 1 256 1 1 0 257
0
0 0 4720 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
4441 0 0
0
0
AAAAABACADAEAFAGAHAIAJAKALAMANAOAPBABBBCBDBEBFBGBHBIBJBKBLBMBNBOBPCACBCCCDCECFCG
CHCICJCKCLCMCNCOCPDADBDCDDDEDFDGDHDIDJDKDLDMDNDODPEAEBECEDEEEFEGEHEIEJEKELEMENEO
EPFAFBFCFDFEFFFGFHFIFJFKFLFMFNFOFPGAGBGCGDGEGFGGGHGIGJGKGLGMGNGOGPHAHBHCHDHEHFHG
HHHIHJHKHLHMHNHOHPIAIBICIDIEIFIGIHIIIJIKILIMINIOIPJAJBJCJDJEJFJGJHJIJJJKJLJMJNJO
JPKAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPLALBLCLDLELFLGLHLILJLKLLLMLNLOLPMAMBMCMDMEMFMG
MHMIMJMKMLMMMNMOMPNANBNCNDNENFNGNHNINJNKNLNMNNNONPOAOBOCODOEOFOGOHOIOJOKOLOMONOO
OPPAPBPCPDPEPFPGPHPIPJPKPLPMPNPOPP
2 +V
167 238 39 0 1 3
0 4
0
0 0 54256 0
4 5.12
-14 -22 14 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
7 Ground~
168 239 153 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
5 SAVE-
218 259 74 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
5 SAVE1
-11 -36 24 -28
0
0
14 *TRAN 0 580m 0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
5394 0 0
0
0
11
11 0 3 0 0 4224 0 1 0 0 0 2
204 74
288 74
9 1 2 0 0 8320 0 1 4 0 0 3
204 101
239 101
239 147
10 1 4 0 0 8320 0 1 3 0 0 3
204 92
238 92
238 48
8 8 5 0 0 4224 0 1 2 0 0 2
138 119
83 119
7 7 6 0 0 4224 0 2 1 0 0 2
83 110
138 110
6 6 7 0 0 4224 0 1 2 0 0 2
138 101
83 101
5 5 8 0 0 4224 0 2 1 0 0 2
83 92
138 92
4 4 9 0 0 4224 0 1 2 0 0 2
138 83
83 83
3 3 10 0 0 4224 0 2 1 0 0 2
83 74
138 74
2 2 11 0 0 4224 0 2 1 0 0 2
83 65
138 65
1 1 12 0 0 4224 0 2 1 0 0 2
83 56
138 56
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 3e-005 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
692 8550464 100 100 0 0
77 66 767 186
0 319 800 572
767 66
77 66
767 126
767 126
0 0
3e-005 0 0 0 3e-005 3e-005
13425 0
2 5e-006 10
6
223 74
0 3 0 -59 1	0 1 0 0
97 119
0 5 0 -39 1	0 4 0 0
102 110
0 6 0 -19 1	0 5 0 0
104 101
0 7 0 4 1	0 6 0 0
108 92
0 8 0 23 1	0 7 0 0
113 83
0 9 0 42 1	0 8 0 0
0 0 100 100 0 0
77 66 767 186
0 0 0 0
767 66
77 66
767 66
767 186
0 0
0.0002 0 0 0 0.0002 0.0002
13425 0
0 5e-005 5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
