CircuitMaker Text
5.6
Probes: 2
V1_1
Transient Analysis
0 186 110 65280
T1_4
Transient Analysis
1 348 110 65535
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
231 152 911 669
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
2 4 0.500000 0.500000
231 411 911 669
12058626 0
0
6 Title:
5 Name:
0
0
0
5
5 xfmr~
219 283 129 0 4 9
0 5 2 2 3
0
0 0 4944 0
7 DEFAULT
-22 -36 27 -28
2 T1
-4 -46 10 -38
0
0
17 %D %1 %2 %3 %4 %S
0
40 alias:XXFMR {PRIT=10 SECT=100 FRAC=TRUE}
0
9

0 1 2 3 4 1 2 3 4 0
88 0 0 0 1 0 0 0
1 T
6641 0 0
2
36626.6 0
0
7 Ground~
168 286 211 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6144 0 0
2
36626.6 1
0
11 Signal Gen~
195 143 116 0 19 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4208 0 0
2
36626.6 2
0
9 Resistor~
219 218 111 0 2 5
0 4 5
0
0 0 880 0
2 1m
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3644 0 0
2
36626.6 3
0
9 Resistor~
219 389 111 0 4 5
0 3 2 0 -1
0
0 0 880 0
3 100
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8720 0 0
2
36626.6 4
0
7
1 0 2 0 0 4096 0 2 0 0 5 2
286 205
286 190
2 0 2 0 0 8192 0 1 0 0 5 3
259 147
249 147
249 190
3 0 2 0 0 0 0 1 0 0 5 3
313 147
318 147
318 190
4 1 3 0 0 4224 0 1 5 0 0 2
313 111
371 111
2 2 2 0 0 12416 0 3 5 0 0 6
174 121
181 121
181 190
415 190
415 111
407 111
1 1 4 0 0 4224 0 4 3 0 0 2
200 111
174 111
1 2 5 0 0 4224 0 1 4 0 0 2
259 111
236 111
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
3900 8550464 100 100 0 0
77 66 977 246
0 403 1024 740
977 66
77 66
977 66
977 246
0 0
4.94359e-315 0 5.4086e-315 1.60186e-314 4.94359e-315 4.94359e-315
12401 0
4 0.001 5
2
187 111
0 4 0 0 1	0 6 0 0
348 111
0 3 0 0 1	0 4 0 0
3420 8550464 100 100 0 0
77 66 977 246
0 403 1024 740
977 66
77 66
977 66
977 246
0 0
0 0 0 0 0 0
12401 0
4 0.001 5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
