CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 480
7 5.000 V
7 5.000 V
3 GND
0 66 640 480
168820736 0
0
0
0
0
0
0
24
10 Ascii Key~
169 47 70 0 11 64
0 7 6 5 4 103 104 105 8 0
0 50
0
0 0 20528 0
0
0
0
0
0
0
0
0
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 -1610612616
0 0 0 512 1 0 0 0
0
8953 0 0
0
0
7 Pulser~
4 243 286 0 12 64
0 10 106 107 9 0 0 32 8 -1
7 1 -1373
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612511
0 0 0 512 1 0 0 0
0
4441 0 0
0
0
8 Hex Key~
166 143 167 0 11 64
0 11 12 13 14 0 0 0 0 0
2 50
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612511
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
8 Hex Key~
166 108 167 0 11 64
0 15 16 17 18 0 0 0 0 0
4 52
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612511
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
8 Hex Key~
166 72 166 0 11 64
0 20 21 22 19 0 0 0 0 0
7 55
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612616
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
8 Hex Key~
166 36 166 0 11 64
0 26 25 24 23 0 0 0 0 0
1 49
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612616
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
8 Hex Key~
166 454 53 0 11 64
0 31 32 33 34 0 0 0 0 0
0 48
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612616
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
8 Hex Key~
166 418 53 0 11 64
0 35 36 37 38 0 0 0 0 0
2 50
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612616
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
5 Delay
94 508 112 0 11 64
0 38 37 36 35 34 33 32 31 30
29 9
5 Delay
1 0 4240 0
0
0
0
0
0
0
0
0
23

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 -1610612712
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
7 Ground~
168 316 287 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -1610612487
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
8 Hex Key~
166 168 52 0 11 64
0 40 41 42 43 0 0 0 0 0
0 48
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612616
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
8 Hex Key~
166 131 52 0 11 64
0 44 45 46 47 0 0 0 0 0
1 49
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612616
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
5 Delay
94 221 113 0 11 64
0 47 46 45 44 43 42 41 40 28
39 9
5 Delay
2 0 4240 0
0
0
0
0
0
0
0
0
23

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 -1610612632
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
14 Logic Display~
6 385 44 0 1 64
10 28
0
0 0 53280 0
0
0
0
0
0
0
0
0
3

0 1 1 -1610612487
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
9 Inverter~
13 451 239 0 2 64
0 27 48
0
0 0 112 90
4 7404
-11 -28 17 -20
0
0
13 VCC=14;GND=7;
11 %D %1 %2 %S
0
0
5 DIP14
64

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0
88 0 0 0 6 1 1 0
1 U
7668 0 0
0
0
6 74LS74
17 509 222 0 12 64
0 132 133 48 28 134 135 136 137 138
29 139 140
0
0 0 4272 0
6 74LS74
-21 -61 21 -53
0
0
13 VCC=14;GND=7;
0
0
0
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 -1610612632
0 0 0 512 1 0 0 0
1 U
4718 0 0
0
0
14 NO PushButton~
191 351 132 0 2 64
0 39 2
0
0 0 20592 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 -1610612495
0 0 0 0 1 0 0 0
1 S
3874 0 0
0
0
14 NO PushButton~
191 299 132 0 2 64
0 2 9
0
0 0 20592 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 -1610612495
0 0 0 0 1 0 0 0
1 S
6671 0 0
0
0
7 Window~
179 362 225 0 11 64
0 27 28 141 142 0 0 0 0 0
0 1
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612632
0 0 0 512 1 0 0 0
0
3789 0 0
0
0
7 Ground~
168 572 286 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -1610612487
0 0 0 0 1 0 0 0
0
4871 0 0
0
0
13 Piezo Buzzer~
174 572 234 0 2 64
10 30 2
0
0 0 20528 270
0
0
0
0
0
0
0
0
5

0 1 2 1 2 -1610612495
0 0 0 0 1 0 0 0
0
3750 0 0
0
0
7 Window~
179 222 223 0 11 64
0 27 28 143 144 0 0 0 0 0
0 1
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612632
0 0 0 512 1 0 0 0
0
8778 0 0
0
0
4 Lock
94 110 236 0 22 64
0 19 22 21 20 18 17 16 15 14
13 12 11 8 7 6 5 4 10 26
25 24 23
4 Lock
3 0 4240 782
0
0
0
0
0
0
0
0
45

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612655
0 0 0 0 1 0 0 0
0
538 0 0
0
0
9 Resistor~
219 498 273 0 4 64
0 27 2 0 -1
9 Resistor~
0 0 4208 0
2 1k
-7 -14 7 -6
0
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -1610612495
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
62
17 4 4 0 0 4288 0 23 0 0 11 2
126 270
126 299
16 3 5 0 0 4288 0 23 0 0 11 2
135 270
135 299
15 2 6 0 0 4288 0 23 0 0 11 2
144 270
144 299
14 1 7 0 0 4288 0 23 0 0 11 2
153 270
153 299
13 5 8 0 0 4288 0 23 0 0 11 2
162 270
162 299
8 5 8 0 0 64 0 1 0 0 11 2
26 94
26 117
4 4 4 0 0 64 0 1 0 0 11 2
50 94
50 117
3 3 5 0 0 64 0 1 0 0 11 2
56 94
56 117
2 2 6 0 0 64 0 1 0 0 11 2
62 94
62 117
1 1 7 0 0 64 0 1 0 0 11 2
68 94
68 117
1 0 1 0 0 8352 0 0 0 0 0 4
77 117
11 117
11 299
179 299
0 4 9 0 0 4096 0 0 2 34 0 3
297 163
297 286
273 286
18 1 10 0 0 8320 0 23 2 0 0 3
108 270
108 277
219 277
1 12 11 0 0 12416 0 3 23 0 0 4
152 191
152 193
162 193
162 206
2 11 12 0 0 12416 0 3 23 0 0 4
146 191
146 197
153 197
153 206
3 10 13 0 0 4224 0 3 23 0 0 4
140 191
140 201
144 201
144 206
4 9 14 0 0 8320 0 3 23 0 0 3
134 191
135 191
135 206
1 8 15 0 0 12416 0 4 23 0 0 4
117 191
117 196
126 196
126 206
2 7 16 0 0 8320 0 4 23 0 0 5
111 191
110 191
110 199
117 199
117 206
3 6 17 0 0 4224 0 4 23 0 0 4
105 191
105 201
108 201
108 206
5 4 18 0 0 4224 0 23 4 0 0 2
99 206
99 191
1 4 19 0 0 4224 0 23 5 0 0 2
63 206
63 190
1 4 20 0 0 12416 0 5 23 0 0 4
81 190
81 196
90 196
90 206
2 3 21 0 0 8320 0 5 23 0 0 5
75 190
76 190
76 200
81 200
81 206
3 2 22 0 0 4224 0 5 23 0 0 4
69 190
69 200
72 200
72 206
22 4 23 0 0 12416 0 23 6 0 0 4
63 270
63 289
27 289
27 190
3 21 24 0 0 4224 0 6 23 0 0 4
33 190
33 284
72 284
72 270
20 2 25 0 0 12416 0 23 6 0 0 4
81 270
81 279
39 279
39 190
1 19 26 0 0 4224 0 6 23 0 0 4
45 190
45 274
90 274
90 270
1 1 27 0 0 12416 0 22 24 0 0 4
268 241
279 241
279 273
480 273
2 0 2 0 0 4096 0 24 0 0 32 2
516 273
558 273
2 1 2 0 0 0 0 21 20 0 0 6
572 265
572 273
558 273
558 273
572 273
572 280
1 0 28 0 0 4096 0 14 0 0 51 2
385 62
385 171
0 11 9 0 0 8320 0 0 9 49 0 5
272 140
272 163
560 163
560 139
546 139
10 10 29 0 0 8320 0 9 16 0 0 5
546 148
552 148
552 203
547 203
547 204
9 1 30 0 0 8320 0 9 21 0 0 3
540 94
572 94
572 203
8 1 31 0 0 8320 0 9 7 0 0 3
476 148
463 148
463 77
2 7 32 0 0 4224 0 7 9 0 0 3
457 77
457 139
476 139
3 6 33 0 0 4224 0 7 9 0 0 3
451 77
451 130
476 130
5 4 34 0 0 8320 0 9 7 0 0 3
476 121
445 121
445 77
1 4 35 0 0 8320 0 8 9 0 0 3
427 77
427 112
476 112
2 3 36 0 0 8320 0 8 9 0 0 3
421 77
421 103
476 103
3 2 37 0 0 8320 0 8 9 0 0 3
415 77
415 94
476 94
1 4 38 0 0 4224 0 9 8 0 0 3
476 85
409 85
409 77
4 0 28 0 0 0 0 16 0 0 51 2
471 213
417 213
1 1 2 0 0 4224 0 18 10 0 0 2
316 140
316 281
2 1 2 0 0 0 0 17 18 0 0 2
334 140
316 140
10 1 39 0 0 4224 0 13 17 0 0 4
259 149
379 149
379 140
368 140
11 2 9 0 0 0 0 13 18 0 0 2
259 140
282 140
2 0 28 0 0 0 0 22 0 0 51 3
268 232
278 232
278 171
2 9 28 0 0 12416 0 19 13 0 0 6
408 234
417 234
417 171
264 171
264 95
253 95
8 1 40 0 0 8320 0 13 11 0 0 3
189 149
177 149
177 76
2 7 41 0 0 4224 0 11 13 0 0 3
171 76
171 140
189 140
3 6 42 0 0 4224 0 11 13 0 0 3
165 76
165 131
189 131
5 4 43 0 0 8320 0 13 11 0 0 3
189 122
159 122
159 76
1 4 44 0 0 8320 0 12 13 0 0 3
140 76
140 113
189 113
2 3 45 0 0 8320 0 12 13 0 0 3
134 76
134 104
189 104
3 2 46 0 0 8320 0 12 13 0 0 3
128 76
128 95
189 95
1 4 47 0 0 4224 0 13 12 0 0 3
189 86
122 86
122 76
2 3 48 0 0 4224 0 15 16 0 0 3
454 221
454 204
471 204
1 0 27 0 0 0 0 15 0 0 30 2
454 257
454 273
1 0 27 0 0 0 0 19 0 0 30 3
408 243
418 243
418 273
7
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 12
273 72 340 122
277 76 330 114
12 Reset
Alarm
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 13
326 72 393 122
330 76 383 114
13 Enable
Alarm
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 5
324 36 383 63
328 40 373 59
5 Armed
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 18
195 22 284 72
199 26 274 64
18 Exit Delay 
Time
-16 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 19
478 25 577 75
482 29 567 67
19 Entry Delay 
Time
-17 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 15
20 116 158 143
24 120 148 139
15 Set Combination
-17 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 18
5 0 129 50
9 4 119 42
18 Input
Combination
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
