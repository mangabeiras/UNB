CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 442 429
7 5.000 V
7 5.000 V
3 GND
0 66 442 429
12058624 0
0
0
0
0
0
0
13
5 SAVE-
218 193 143 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
25 *Combine
*TRAN -13m 6.62
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 95 145 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
25 *Combine
*TRAN -13m 6.62
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
2 +V
167 142 239 0 1 3
0 10
0
0 0 54112 -19276
4 -15V
-12 0 16 8
2 V1
-7 12 7 20
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3618 0 0
0
0
2 +V
167 21 160 0 1 3
0 11
0
0 0 54112 7168
3 -8V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6153 0 0
0
0
2 +V
167 291 32 0 1 3
0 6
0
0 0 54112 0
2 6V
15 -2 29 6
2 V3
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
2 +V
167 142 143 0 1 3
0 9
0
0 0 54112 0
3 15V
-11 -13 10 -5
2 V4
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7734 0 0
0
0
7 Ground~
168 93 237 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
8 Op-Amp7~
219 142 187 0 7 15
0 2 8 9 10 3 4 5
8 Op-Amp7~
0 0 832 0
6 LM301A
6 -24 48 -16
2 U1
20 -34 34 -26
0
0
26 %D %1 %2 %3 %4 %5 %6 %7 %S
0
0
4 DIP8
15

0 3 2 7 4 6 1 8 3 2
7 4 6 1 8 -33686019
88 0 0 256 1 1 0 0
1 U
3747 0 0
0
0
10 Capacitor~
219 144 105 0 2 5
0 8 3
10 Capacitor~
0 0 832 0
5 .05uF
-19 -18 16 -10
2 C1
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
3549 0 0
0
0
10 Capacitor~
219 187 226 0 2 5
0 5 4
10 Capacitor~
0 0 832 0
5 4.7pF
-16 10 19 18
2 C2
-6 -18 8 -10
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
7931 0 0
0
0
4 PUT~
219 143 62 0 3 64
0 3 7 8
4 PUT~
0 0 832 26894
6 2N6027
-17 -23 25 -15
4 PUT1
-8 -35 20 -27
0
0
14 %D %1 %2 %3 %S
0
0
8 TO-226AA
4

0 1 2 3 0
88 0 0 0 1 0 0 0
3 PUT
9325 0 0
0
0
9 Resistor~
219 61 181 0 3 5
0 11 8 1
9 Resistor~
0 0 4960 0
2 5k
-7 -12 7 -4
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 229 52 0 4 5
0 7 6 0 1
9 Resistor~
0 0 4960 0
2 5k
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3834 0 0
0
0
13
2 0 3 0 0 4096 0 9 0 0 2 2
153 105
193 105
5 1 3 0 0 8320 0 8 11 0 0 4
160 187
193 187
193 62
157 62
6 2 4 0 0 4224 0 8 10 0 0 4
158 179
206 179
206 226
196 226
7 1 5 0 0 8320 0 8 10 0 0 4
158 195
172 195
172 226
178 226
2 1 6 0 0 4224 0 13 5 0 0 3
247 52
291 52
291 41
2 1 7 0 0 4224 0 11 13 0 0 2
157 52
211 52
1 0 8 0 0 4096 0 9 0 0 8 2
135 105
95 105
3 0 8 0 0 8320 0 11 0 0 12 3
129 62
95 62
95 181
3 1 9 0 0 4224 0 8 6 0 0 2
142 174
142 152
4 1 10 0 0 4224 0 8 3 0 0 2
142 200
142 224
1 1 2 0 0 8320 0 8 7 0 0 3
124 193
93 193
93 231
2 2 8 0 0 0 0 12 8 0 0 2
79 181
124 181
1 1 11 0 0 8320 0 4 12 0 0 3
21 169
21 181
43 181
0
0
16 2 0
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 0.0005 5e-005 5e-005 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
3904 8550464 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
4.80864e-315 0 5.4086e-315 0 4.80864e-315 5.4086e-315
16 0
4 0.0001 10
1
175 52
0 7 0 0 1	0 6 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
