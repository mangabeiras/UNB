CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 640 413
7 5.000 V
7 5.000 V
3 GND
2500 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 413
12058634 0
0
0
0
0
0
0
25
5 SAVE-
218 416 134 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
10 *TRAN 6 12
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
7 Ground~
168 103 247 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
11 Signal Gen~
195 48 217 0 19 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 -1090519040 1050253722
20
1 1000 -0.5 0.3 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 320 0
12 -800m/-200mV
-41 -28 43 -20
2 V1
-7 -38 7 -30
0
0
43 %D %1 %2 DC 0 SIN(-500m 300m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
11 Signal Gen~
195 48 155 0 19 64
0 13 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1203982336 0 1056964608
20
1 100000 0 0.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 320 0
11 -500m/500mV
-38 -28 39 -20
2 V2
-7 -38 7 -30
0
0
41 %D %1 %2 DC 0 SIN(0 500m 100k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
7 Ground~
168 416 231 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
7 Ground~
168 281 106 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
7 Ground~
168 158 67 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
7 Ground~
168 273 252 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
2 +V
167 391 298 0 1 64
0 9
0
0 0 53600 -19276
3 -8V
7 -10 28 -2
2 V3
10 -20 24 -12
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
2 +V
167 442 23 0 1 64
0 16
0
0 0 53600 0
4 +12V
8 -3 36 5
2 V4
15 -13 29 -5
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
10 Capacitor~
219 122 150 0 2 64
0 13 11
10 Capacitor~
0 0 320 0
4 .1uF
-15 -19 13 -11
2 C1
-8 -29 6 -21
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
9325 0 0
0
0
10 Capacitor~
219 281 74 0 2 64
0 12 2
10 Capacitor~
0 0 320 26894
4 .1uF
14 -3 42 5
2 C2
21 -13 35 -5
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
8903 0 0
0
0
13 Var Resistor~
219 181 239 0 3 64
0 14 9 15
13 Var Resistor~
0 0 320 -19276
7 50k 80%
-24 -20 25 -12
2 R1
-7 -30 7 -22
0
0
32 %DA %1 %2 40000
%DB %2 %3 10000
0
0
4 SIP3
7

0 1 2 3 1 2 3 -33686019
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
6 MC1496
219 345 150 0 10 64
0 4 12 11 3 10 9 8 7 6
5
6 MC1496
0 0 12480 0
6 MC1496
-21 -42 21 -34
2 U1
-7 -52 7 -44
0
0
36 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %10 %S
0
0
5 DIP14
21

0 2 8 10 1 4 14 5 12 6
3 2 8 10 1 4 14 5 12 6
3 -33686019
88 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
9 Resistor~
219 198 46 0 3 64
0 2 12 -1
9 Resistor~
0 0 352 0
2 1k
-7 -12 7 -4
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 214 108 0 2 64
0 11 12
9 Resistor~
0 0 352 0
2 51
-7 -12 7 -4
2 R3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 342 46 0 4 64
0 12 16 0 1
9 Resistor~
0 0 352 0
2 1k
-7 -12 7 -4
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 343 102 0 2 64
0 4 5
9 Resistor~
0 0 352 0
2 1k
-7 -12 7 -4
2 R5
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 416 79 0 4 64
0 6 16 0 1
9 Resistor~
0 0 352 90
4 3.9k
6 -5 34 3
2 R6
13 -15 27 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 470 79 0 4 64
0 7 16 0 1
9 Resistor~
0 0 352 90
4 3.9k
7 -5 35 3
2 R7
13 -17 27 -9
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 416 192 0 3 64
0 2 8 -1
9 Resistor~
0 0 352 90
4 6.8k
6 -2 34 6
2 R8
12 -12 26 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 296 200 0 3 64
0 2 10 -1
9 Resistor~
0 0 352 90
2 51
7 -5 21 3
2 R9
7 -15 21 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 246 200 0 3 64
0 2 3 -1
9 Resistor~
0 0 352 90
2 51
6 -5 20 3
3 R10
3 -15 24 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 209 197 0 2 64
0 14 10
9 Resistor~
0 0 352 90
3 750
6 -1 27 7
3 R11
6 -12 27 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 152 198 0 2 64
0 15 3
9 Resistor~
0 0 352 90
3 750
6 -2 27 6
3 R12
4 -11 25 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
31
1 0 2 0 0 4096 0 8 0 0 21 2
273 246
273 231
1 0 3 0 0 4096 0 3 0 0 12 4
79 212
140 212
140 159
152 159
2 0 2 0 0 4096 0 3 0 0 4 2
79 222
103 222
1 2 2 0 0 4224 0 2 4 0 0 3
103 241
103 160
79 160
1 1 4 0 0 8320 0 14 18 0 0 4
313 132
305 132
305 102
325 102
10 2 5 0 0 8320 0 14 18 0 0 4
377 132
385 132
385 102
361 102
9 1 6 0 0 8320 0 14 19 0 0 3
377 141
416 141
416 97
8 1 7 0 0 4224 0 14 20 0 0 3
377 150
470 150
470 97
7 2 8 0 0 4224 0 14 21 0 0 3
377 159
416 159
416 174
6 1 9 0 0 8192 0 14 9 0 0 3
377 168
391 168
391 283
5 2 10 0 0 4224 0 14 24 0 0 3
313 168
209 168
209 179
4 2 3 0 0 4224 0 14 25 0 0 3
313 159
152 159
152 180
3 2 11 0 0 4224 0 14 11 0 0 2
313 150
131 150
2 0 12 0 0 8192 0 14 0 0 30 3
313 141
246 141
246 46
1 1 13 0 0 4224 0 4 11 0 0 2
79 150
113 150
2 0 10 0 0 0 0 22 0 0 11 2
296 182
296 168
2 0 3 0 0 0 0 23 0 0 12 2
246 182
246 159
2 0 9 0 0 8320 0 13 0 0 10 3
183 243
183 273
391 273
1 1 14 0 0 4224 0 24 13 0 0 3
209 215
209 231
199 231
1 3 15 0 0 4224 0 25 13 0 0 3
152 216
152 231
163 231
1 1 2 0 0 0 0 23 22 0 0 4
246 218
246 231
296 231
296 218
1 1 2 0 0 0 0 21 5 0 0 2
416 210
416 225
1 0 11 0 0 0 0 16 0 0 13 3
196 108
182 108
182 150
2 0 12 0 0 0 0 16 0 0 14 2
232 108
246 108
2 1 2 0 0 0 0 12 6 0 0 2
281 83
281 100
1 0 12 0 0 0 0 12 0 0 30 2
281 65
281 46
1 0 16 0 0 4096 0 10 0 0 29 2
442 32
442 46
2 0 16 0 0 4096 0 19 0 0 29 2
416 61
416 46
2 2 16 0 0 4224 0 17 20 0 0 3
360 46
470 46
470 61
2 1 12 0 0 4224 0 15 17 0 0 2
216 46
324 46
1 1 2 0 0 0 0 15 7 0 0 3
180 46
158 46
158 61
1
-16 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
14 24 144 53
18 28 138 47
12 AM Modulator
0
17 0 1
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 0.002 2e-006 2e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
