CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 325 452
8  5.000 V
8  5.000 V
3 GND
125 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 325 452
9961490 0
0
0
0
0
0
0
9
5 SAVE-
218 246 77 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
24 *Combine
*TRAN -168 169
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 105 72 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
24 *Combine
*TRAN -168 169
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
7 Ground~
168 171 184 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
11 Signal Gen~
195 64 99 0 19 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1114636288 0 1126825984
20
1 60 0 170 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
9 -170/170V
-31 -28 32 -20
2 V1
-7 -38 7 -30
0
0
38 %D %1 %2 DC 0 SIN(0 170 60 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
4 SCR~
219 245 107 0 3 7
0 5 4 2
4 SCR~
0 0 832 0
6 2N5064
12 0 54 8
4 SCR1
19 -10 47 -2
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
88 0 0 256 1 1 0 0
3 SCR
5394 0 0
0
0
13 Var Resistor~
219 166 69 0 3 7
0 3 3 5
13 Var Resistor~
0 0 832 90
8 100k 40%
8 -4 64 4
2 R1
29 -14 43 -6
0
0
32 %DA %1 %2 40000
%DB %2 %3 60000
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
10 Polar Cap~
219 172 140 0 2 5
0 3 2
10 Polar Cap~
0 0 832 270
5 .25uF
10 4 45 12
2 C1
21 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
9914 0 0
0
0
6 Diode~
219 207 113 0 2 5
0 3 4
6 Diode~
0 0 832 0
6 1N4934
-20 -18 22 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 0 0 0 1 1 0 0
1 D
3747 0 0
0
0
9 Resistor~
219 137 35 0 2 5
0 6 5
9 Resistor~
0 0 4960 0
3 100
-10 -12 11 -4
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3549 0 0
0
0
10
0 2 3 0 0 8320 0 0 6 3 0 4
171 113
140 113
140 67
160 67
2 2 4 0 0 4224 0 8 5 0 0 2
217 113
232 113
1 0 3 0 0 0 0 8 0 0 5 2
197 113
171 113
3 0 5 0 0 4096 0 6 0 0 9 2
170 47
170 35
1 1 3 0 0 0 0 7 6 0 0 4
171 130
171 85
170 85
170 83
2 0 2 0 0 4096 0 7 0 0 8 2
171 147
171 161
1 0 2 0 0 4096 0 3 0 0 8 2
171 178
171 161
3 2 2 0 0 8320 0 5 4 0 0 5
245 119
245 161
104 161
104 104
95 104
2 1 5 0 0 4224 0 9 5 0 0 3
155 35
245 35
245 95
1 1 6 0 0 8320 0 4 9 0 0 4
95 94
104 94
104 35
119 35
0
0
16 0 0
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 0.04 0.001 0.001
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2188 8526400 100 100 0 0
98 66 278 156
325 66 640 291
278 66
98 66
278 66
278 156
0 0
5.06792e-315 0 5.30499e-315 1.58155e-314 5.06792e-315 5.06792e-315
8313 0
4 0.01 100
1
155 35
0 5 0 0 1	0 9 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
