CircuitMaker Text
5.6
Probes: 3
Signal
Transient Analysis
0 118 58 65280
LED1
Transient Analysis
1 557 117 65535
LED2
Transient Analysis
2 450 102 16776960
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 9 100 10
231 152 911 669
7 5.000 V
7 5.000 V
3 GND
1.66667 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
2 4 0.500000 0.500000
231 411 911 669
11010066 0
0
0
0
0
0
0
15
12 NPN Trans:C~
219 226 57 0 3 7
0 8 10 7
12 NPN Trans:C~
0 0 848 0
6 2N3904
20 -4 62 4
2 Q1
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
3577 0 0
2
36626.5 10
0
4 LED~
171 455 140 0 2 5
10 4 9
0
0 0 624 0
4 LED2
10 -16 38 -8
2 D2
9 -18 23 -10
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3727 0 0
2
36626.5 9
0
4 LED~
171 556 142 0 2 5
12 5 9
0
0 0 624 0
4 LED2
10 -16 38 -8
2 D1
8 -18 22 -10
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4144 0 0
2
36626.5 8
0
7 Ground~
168 218 173 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4788 0 0
2
36626.5 7
0
2 +V
167 231 25 0 1 3
0 8
0
0 0 53616 0
3 +5V
12 -2 33 6
2 V2
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
359 0 0
2
36626.5 6
0
7 Ground~
168 101 79 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
842 0 0
2
36626.5 5
0
12 SPST Switch~
165 351 121 0 2 11
0 6 4
0
0 0 20592 512
0
2 S1
-7 -28 7 -20
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6593 0 0
2
36626.5 4
0
4 .IC~
207 258 104 0 1 3
0 6
0
0 0 53584 0
2 0V
-7 -15 7 -7
4 CMD1
-14 -25 14 -17
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
3 CMD
4896 0 0
2
36626.5 3
0
9 2-In NOR~
219 314 93 0 3 21
0 7 6 5
0
0 0 112 0
6 74LS02
-21 -24 21 -16
3 U1A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 1 0
1 U
3822 0 0
2
36626.5 2
0
9 2-In NOR~
219 407 102 0 3 21
0 5 5 4
0
0 0 112 0
6 74LS02
-21 -24 21 -16
3 U1B
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
5367 0 0
2
36626.5 1
0
11 Signal Gen~
195 54 62 0 64 64
0 3 2 1 86 -8 8 0 0 0
0 0 0 0 0 0 0 1065353216 0 1083179008
1056964608 1020054733 1020054733 1045220557 1065353216 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 264
20
0 1 0 4.5 0.5 0.025 0.025 0.2 1 0
0 0 0 0 0 0 0 0 0 0
0
0 0 336 0
6 0/4.5V
-20 -28 22 -20
2 V1
-7 -38 7 -30
0
0
46 %D %1 %2 DC 0 PULSE(0 4.5 500m 25m 25m 200m 1)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6131 0 0
2
36626.5 0
0
9 Resistor~
219 176 57 0 2 11
0 3 10
9 Resistor~
0 0 880 0
2 1k
-7 -12 7 -4
2 R4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
3114 0 0
2
36626.5 14
0
9 Resistor~
219 231 141 0 3 11
0 2 7 -1
9 Resistor~
0 0 880 90
3 470
7 1 28 9
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
7771 0 0
2
36626.5 13
0
9 Resistor~
219 280 145 0 3 11
0 2 6 -1
9 Resistor~
0 0 880 90
3 470
4 3 25 11
2 R2
6 -7 20 1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
7563 0 0
2
36626.5 12
0
9 Resistor~
219 412 166 0 3 11
0 2 9 -1
9 Resistor~
0 0 880 0
3 150
-10 -12 11 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
9849 0 0
2
36626.5 11
0
19
2 1 2 0 0 4112 0 11 6 0 0 3
85 67
101 67
101 73
1 1 3 0 0 4240 0 12 11 0 0 2
158 57
85 57
3 1 4 0 0 8208 0 10 2 0 0 3
446 102
455 102
455 130
1 2 5 0 0 4112 0 10 10 0 0 4
394 93
373 93
373 111
394 111
3 0 5 0 0 16 0 9 0 0 4 2
353 93
373 93
2 2 6 0 0 8208 0 9 14 0 0 3
301 102
280 102
280 127
1 0 7 0 0 4240 0 9 0 0 18 2
301 84
231 84
1 0 2 0 0 16 0 4 0 0 17 3
218 167
218 166
231 166
1 0 6 0 0 16 0 8 0 0 6 3
258 116
258 121
280 121
1 0 5 0 0 8336 0 3 0 0 5 4
556 132
556 56
373 56
373 93
1 0 6 0 0 4240 0 7 0 0 6 2
334 121
280 121
2 0 4 0 0 4240 0 7 0 0 3 2
368 121
455 121
1 1 8 0 0 4240 0 5 1 0 0 2
231 34
231 39
2 0 9 0 0 4112 0 2 0 0 15 2
455 150
455 166
2 2 9 0 0 4240 0 15 3 0 0 3
430 166
556 166
556 152
1 0 2 0 0 16 0 14 0 0 17 2
280 163
280 166
1 1 2 0 0 8336 0 13 15 0 0 3
231 159
231 166
394 166
3 2 7 0 0 16 0 1 13 0 0 2
231 75
231 123
2 2 10 0 0 4240 0 12 1 0 0 2
194 57
208 57
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 6
99 41 150 57
99 41 150 57
6 Signal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 4
455 97 490 113
455 97 490 113
4 LED2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 4
556 82 591 98
556 82 591 98
4 LED1
-11 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
121 58 191 78
125 62 188 76
9 Probe Tip
-20 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 11
371 19 512 54
375 23 507 50
11 Logic Probe
19 .OPTIONS TRTOL=10

16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 3 0.025 0.025
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
164 8526400 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 89
617 98
0 0
0 0 0 0 0 0
13433 0
2 0.5 5
3
109 128
0 3 0 16 1	0 14 0 0
482 168
0 5 0 0 1	0 20 0 0
431 173
0 4 0 -15 1	0 13 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
