CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 100 3
0 70 640 452
7 5.000 V
7 5.000 V
3 GND
0 70 640 452
143654914 0
0
0
0
0
0
0
5
9 CA 7-Seg~
184 215 109 1 18 19
10 8 7 6 5 4 3 2 21 16
0 0 0 0 0 0 0 2 1
0
0 0 20592 0
5 REDCA
16 -41 51 -33
5 DISP1
16 -51 51 -43
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
8953 0 0
0
0
9 CC 7-Seg~
183 383 108 1 18 19
10 15 14 13 12 11 10 9 22 16
1 1 1 1 1 1 1 2 1
0
0 0 20592 0
5 REDCC
16 -41 51 -33
5 DISP2
16 -51 51 -43
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
4441 0 0
0
0
6 74LS48
188 318 208 0 14 29
0 18 17 19 20 23 24 9 10 11
12 13 14 15 25
0
0 0 12512 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -70 7 -62
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 -33686019
65 0 0 512 1 1 0 0
1 U
3618 0 0
0
0
6 74LS47
187 150 205 0 14 29
0 18 17 19 20 26 27 2 3 4
5 6 7 8 28
0
0 0 12512 0
6 74LS47
-21 -60 21 -52
2 U2
-7 -70 7 -62
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 -33686019
65 0 0 512 1 1 0 0
1 U
6153 0 0
0
0
9 Data Seq~
170 41 58 0 17 21
0 29 30 31 16 18 17 19 20 32
33 18 1 20 1 1 0 33
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -54 10 -46
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
0
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 0 0 0 0
2 DS
5394 0 0
0
0
AAAABAABBBACBCADBDAEBEAFBFAGBGAHBHAIBIAJBJAAAAAAAAAAAAAAAAAAAAAAAA
24
7 7 2 0 0 8320 0 1 4 0 0 3
230 145
230 169
188 169
8 6 3 0 0 4224 0 4 1 0 0 3
188 178
224 178
224 145
5 9 4 0 0 4224 0 1 4 0 0 3
218 145
218 187
188 187
10 4 5 0 0 8320 0 4 1 0 0 3
188 196
212 196
212 145
3 11 6 0 0 4224 0 1 4 0 0 3
206 145
206 205
188 205
12 2 7 0 0 8320 0 4 1 0 0 3
188 214
200 214
200 145
13 1 8 0 0 8320 0 4 1 0 0 3
188 223
194 223
194 145
7 7 9 0 0 4224 0 3 2 0 0 3
350 172
398 172
398 144
6 8 10 0 0 8320 0 2 3 0 0 3
392 144
392 181
350 181
9 5 11 0 0 8320 0 3 2 0 0 3
350 190
386 190
386 144
4 10 12 0 0 4224 0 2 3 0 0 3
380 144
380 199
350 199
11 3 13 0 0 8320 0 3 2 0 0 3
350 208
374 208
374 144
2 12 14 0 0 4224 0 2 3 0 0 3
368 144
368 217
350 217
13 1 15 0 0 8320 0 3 2 0 0 3
350 226
362 226
362 144
0 9 16 0 0 4096 0 0 1 16 0 2
215 58
215 73
4 9 16 0 0 4224 0 5 2 0 0 3
73 58
383 58
383 66
6 2 17 0 0 8192 0 5 4 0 0 4
73 76
92 76
92 178
118 178
1 0 18 0 0 12416 0 3 0 0 22 5
286 172
253 172
253 263
86 263
86 169
0 2 17 0 0 8320 0 0 3 17 0 5
92 178
92 268
259 268
259 181
286 181
3 0 19 0 0 12416 0 3 0 0 23 5
286 190
266 190
266 273
99 273
99 187
0 4 20 0 0 8320 0 0 3 24 0 5
104 196
104 278
272 278
272 199
286 199
1 5 18 0 0 0 0 4 5 0 0 4
118 169
86 169
86 67
73 67
3 7 19 0 0 0 0 4 5 0 0 4
118 187
98 187
98 85
73 85
8 4 20 0 0 0 0 5 4 0 0 4
73 94
104 94
104 196
118 196
0
0
16 0 1
0
0
3 Vin
-1.5 -0.7 0.01
3 Vcc
10 14 1
100 0 1 100000
0 2e-005 8e-008 8e-008 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
3112 8550464 100 100 0 0
77 66 617 126
19 481 659 674
617 66
77 66
617 66
617 126
0 0
0 0 0 0 0 0
16 0
4 5e-006 2
1
194 158
0 8 0 0 2	0 7 0 0
1084 8550464 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 67
617 126
0 0
4.4781e-315 0 5.54867e-315 5.54829e-315 4.4781e-315 5.23039e-315
0 0
4 5e-005 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
