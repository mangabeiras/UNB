CircuitMaker Text
5.6
Probes: 5
V1_1
Operating Point
0 123 63 65280
V3_1
Operating Point
1 151 65 65535
V2_1
Operating Point
2 175 60 16776960
U2_5
Operating Point
3 303 65 16711935
U1_3
Operating Point
4 303 165 11184640
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
245 80 857 634
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
2 4 0.500000 0.500000
245 357 857 634
12058626 0
0
6 Title:
5 Name:
0
0
0
9
10 divider:A~
219 253 74 0 6 13
0 6 5 7 5 3 2
0
0 0 54096 0
6 DIVIDE
-12 -31 30 -23
2 U2
2 -41 16 -33
0
0
41 %D %%vd(%1,%2) %%vd(%3,%4) %%vd(%5,%6) %M
0
12 type:divider
0
13

0 0 0 0 0 0 0 0 0 0
0 0 0 0
65 0 0 0 1 0 0 0
1 U
9132 0 0
2
36626.4 0
0
8 divider~
219 252 164 0 3 7
0 6 7 4
0
0 0 54096 0
6 DIVIDE
-14 -31 28 -23
2 U1
0 -41 14 -33
0
0
14 %D %1 %2 %3 %M
0
12 type:divider
0
7

0 0 0 0 0 0 0 0
65 0 0 0 1 0 0 0
1 U
4186 0 0
2
36626.4 1
0
7 Ground~
168 339 107 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5408 0 0
2
36626.4 2
0
7 Ground~
168 370 204 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8364 0 0
2
36626.4 3
0
2 +V
167 151 40 0 1 3
0 6
0
0 0 54256 0
1 2
-4 -22 3 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7573 0 0
2
36626.4 4
0
2 +V
167 174 42 0 1 3
0 5
0
0 0 54256 0
2 -1
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4139 0 0
2
36626.4 5
0
2 +V
167 123 39 0 1 3
0 7
0
0 0 54256 0
1 4
-4 -22 3 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3911 0 0
2
36626.4 6
0
9 Resistor~
219 335 164 0 4 5
0 4 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7162 0 0
2
36626.4 7
0
9 Resistor~
219 331 65 0 4 5
0 3 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7367 0 0
2
36626.4 8
0
11
1 0 2 0 0 4096 0 3 0 0 3 3
339 101
339 83
338 83
1 2 2 0 0 4096 0 4 8 0 0 3
370 198
370 164
353 164
2 6 2 0 0 12416 0 9 1 0 0 4
349 65
365 65
365 83
291 83
5 1 3 0 0 4224 0 1 9 0 0 2
291 65
313 65
3 1 4 0 0 4224 0 2 8 0 0 2
290 164
317 164
2 0 5 0 0 4224 0 1 0 0 7 2
229 65
174 65
1 4 5 0 0 0 0 6 1 0 0 3
174 51
174 92
229 92
1 0 6 0 0 4096 0 1 0 0 11 2
229 56
151 56
3 0 7 0 0 4096 0 1 0 0 10 2
229 83
123 83
2 1 7 0 0 8320 0 2 7 0 0 3
228 173
123 173
123 48
1 1 6 0 0 8320 0 2 5 0 0 3
228 155
151 155
151 49
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1392 1210432 100 100 0 0
0 0 0 0
1 57 162 127
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 3
1
306 164
0 4 0 0 1	0 5 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
