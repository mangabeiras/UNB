CircuitMaker Text
5.6
Probes: 5
U1_6
DC Sweep
0 303 89 65280
U1_6
Operating Point
0 303 89 65280
U1_6
Transient Analysis
0 303 89 65280
U1_6
Fourier Analysis
0 303 89 65280
out
AC Analysis
0 304 92 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 300 100 10
245 80 925 597
7 5.000 V
7 5.000 V
3 GND
500 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
2 4 0.500000 0.500000
245 339 925 597
9961488 4
0
0
0
0
0
0
12
11 Signal Gen~
195 40 130 0 19 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1036831949
20
1 1000 0 0.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -100m/100mV
-38 -28 39 -20
2 V1
-7 -38 7 -30
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
398 0 0
2
36626.5 0
0
7 Ground~
168 176 179 0 1 3
0 2
0
0 0 49264 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3479 0 0
2
36626.5 2
0
7 Ground~
168 88 161 0 1 3
0 2
0
0 0 49264 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8546 0 0
2
36626.5 3
0
2 +V
167 233 168 0 1 3
0 11
0
0 0 50032 -19276
4 -15V
-13 0 15 8
2 V2
-5 10 9 18
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9272 0 0
2
36626.5 4
0
2 +V
167 233 86 0 1 3
0 10
0
0 0 50032 0
4 +15V
-14 -13 14 -5
2 V3
-5 -23 9 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3206 0 0
2
36626.5 5
0
8 Op-Amp7~
219 233 119 0 7 15
0 4 7 10 11 3 9 8
8 Op-Amp7~
0 0 848 0
6 LM301A
6 -24 48 -16
2 U1
20 -34 34 -26
0
0
26 %D %1 %2 %3 %4 %5 %6 %7 %S
0
0
4 DIP8
15

0 3 2 7 4 6 1 8 3 2
7 4 6 1 8 -33686019
88 0 0 256 1 1 0 0
1 U
3379 0 0
2
36626.5 6
0
10 Capacitor~
219 284 137 0 2 5
0 9 8
10 Capacitor~
0 0 848 26894
4 50pF
12 0 40 8
2 C1
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
3225 0 0
2
36626.5 7
0
10 Capacitor~
219 176 152 0 2 5
0 2 4
10 Capacitor~
0 0 848 90
6 .001uF
7 2 49 10
2 C2
21 -9 35 -1
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 1 0 0
1 C
7574 0 0
2
36626.5 8
0
10 Capacitor~
219 217 29 0 2 5
0 6 3
10 Capacitor~
0 0 848 0
6 .002uF
-22 -18 20 -10
2 C3
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 1 0 0
1 C
731 0 0
2
36626.5 9
0
9 Resistor~
219 254 59 0 2 5
0 7 3
9 Resistor~
0 0 880 0
3 22k
-10 -12 11 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
3749 0 0
2
36626.5 10
0
9 Resistor~
219 99 125 0 2 5
0 5 6
9 Resistor~
0 0 880 0
3 10k
-10 -12 11 -4
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
5242 0 0
2
36626.5 11
0
9 Resistor~
219 151 125 0 2 5
0 6 4
9 Resistor~
0 0 880 0
3 10k
-10 -12 11 -4
2 R3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
3731 0 0
2
36626.5 12
0
14
1 1 2 0 0 4096 0 8 2 0 0 2
176 161
176 173
0 2 4 0 0 4096 0 0 8 8 0 2
176 125
176 143
2 1 2 0 0 8320 0 1 3 0 0 3
71 135
88 135
88 155
1 1 5 0 0 4224 0 11 1 0 0 2
81 125
71 125
1 0 6 0 0 8320 0 9 0 0 7 3
208 29
124 29
124 125
2 0 3 0 0 4096 0 10 0 0 12 2
272 59
303 59
1 2 6 0 0 0 0 12 11 0 0 2
133 125
117 125
1 2 4 0 0 4224 0 6 12 0 0 2
215 125
169 125
1 2 7 0 0 8320 0 10 6 0 0 4
236 59
196 59
196 113
215 113
2 7 8 0 0 8320 0 7 6 0 0 5
284 146
284 149
262 149
262 127
249 127
6 1 9 0 0 4224 0 6 7 0 0 3
249 111
284 111
284 128
5 2 3 0 0 8320 0 6 9 0 0 4
251 119
303 119
303 29
226 29
3 1 10 0 0 4224 0 6 5 0 0 2
233 106
233 95
4 1 11 0 0 4224 0 6 4 0 0 2
233 132
233 153
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 3
303 97 330 113
303 97 330 113
3 out
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 72
341 64 541 128
345 68 537 116
72 Bessel:      C3=.0013uF
Butterworth: C3=.002uF
Chebyshev:   C3=.0068uF
-16 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 23
366 23 516 76
370 27 510 65
23 Low-pass
Active Filter
0
8 0 0
0
0
0
0 0 0
0
0 0 0
60 1 1 1e+07
0 0.01 2.5e-05 2.5e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1656 4397120 100 100 0 0
98 66 616 126
0 259 640 452
615 66
98 66
616 66
616 126
0 0
0 0 0 0 0 0
12403 0
4 3e+06 5e+06
1
303 86
0 6 0 0 2	0 12 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
