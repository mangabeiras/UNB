CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 800 319
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 800 319
9961490 0
0
6 Title:
5 Name:
0
0
0
9
11 Signal Gen~
195 41 98 0 64 64
0 5 2 3 86 -8 8 0 0 0
0 0 0 0 0 0 0 1176256512 0 1065353216
1084227584 1148846080 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
20
0 10000 0 1 5 1000 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
32 %D %1 %2 DC 0 SFFM(0 1 10k 5 1k)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
12 F->V Source~
219 166 94 0 4 9
0 5 2 4 2
0
0 0 592 0
4 FCVS
34 -2 62 6
2 V2
29 0 43 8
0
0
17 %D %1 %2 %3 %4 %S
0
29 alias:XFTOV {VIL=0.1 VIH=0.2}
0
9

0 1 2 3 4 1 2 3 4 0
88 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 155 167 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
5 SAVE-
218 112 59 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
22 *Combine
*TRAN -1 1 0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
4 SAVE
6153 0 0
0
0
5 SAVE-
218 316 59 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
17 *TRAN 9.32 11.3 0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
4 SAVE
5394 0 0
0
0
10 Capacitor~
219 298 99 0 2 5
0 2 3
0
0 0 848 90
2 1u
14 0 28 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
4 .IC~
207 283 31 0 1 3
0 3
0
0 0 54096 0
2 10
-7 -16 7 -8
4 CMD1
-14 -26 14 -18
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
3 CMD
9914 0 0
0
0
9 Resistor~
219 343 105 0 4 5
0 3 2 0 -1
0
0 0 880 270
4 1meg
2 0 30 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 246 60 0 2 5
0 4 3
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
10
1 0 3 0 0 4096 0 7 0 0 3 2
283 43
283 60
1 3 4 0 0 4224 0 9 2 0 0 3
228 60
175 60
175 70
2 1 3 0 0 4224 0 9 8 0 0 3
264 60
343 60
343 87
1 0 2 0 0 4096 0 6 0 0 10 2
298 108
298 137
2 0 3 0 0 0 0 6 0 0 3 2
298 90
298 60
1 0 2 0 0 0 0 3 0 0 10 2
155 161
155 137
4 0 2 0 0 0 0 2 0 0 10 2
175 124
175 137
2 0 2 0 0 0 0 2 0 0 10 2
139 124
139 137
1 1 5 0 0 12416 0 1 2 0 0 5
72 93
85 93
85 59
139 59
139 70
2 2 2 0 0 8320 0 8 1 0 0 5
343 123
343 137
86 137
86 103
72 103
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 1e-006 1e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
3048 8550464 100 100 0 0
77 66 767 186
0 319 800 572
767 66
77 66
767 66
767 186
0 0
0.005 0 15 -3 0.005 0.005
12401 0
4 0.001 10
2
134 59
0 5 0 0 3	0 9 0 0
318 60
0 3 0 0 1	0 3 0 0
2780 8550464 100 100 0 0
77 66 767 186
0 319 800 572
767 66
77 66
767 66
767 186
0 0
0.005 0 15 -3 0.005 0.005
12401 0
4 0.001 10
2
134 59
0 5 0 0 3	0 9 0 0
318 60
0 3 0 0 1	0 3 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
