CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 100 3
0 66 640 452
7 5.000 V
7 5.000 V
3 GND
0 66 640 452
42991616 0
0
0
0
0
0
0
29
7 Ground~
168 427 131 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
14 NO PushButton~
191 56 110 0 2 64
0 6 2
0
0 0 20592 512
0
0
0
0
0
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
1 S
4441 0 0
0
0
6 74LS74
17 56 277 0 12 64
0 30 31 6 8 32 33 34 35 16
36 37 38
0
0 0 4272 0
6 74LS74
-21 -61 21 -53
0
0
13 VCC=14;GND=7;
0
0
0
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 -33686019
0 0 0 512 1 0 0 0
1 U
3618 0 0
0
0
11 2-Input OR~
1 191 78 0 3 64
0 17 8 18
0
0 0 48 512
6 74LS32
-18 -25 24 -17
0
0
13 VCC=14;GND=7;
0
0
0
5 DIP14
64

0 1 2 3 1 2 3 4 5 6
10 9 8 13 12 11 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0
0 0 0 0 4 1 3 0
1 U
6153 0 0
0
0
7 Pulser~
4 288 27 0 10 64
0 39 40 7 41 0 0 5 5 2
7
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -33686019
0 0 0 512 1 0 0 0
0
5394 0 0
0
0
12 2-Input AND~
0 135 59 0 3 64
0 7 18 19
0
0 0 48 512
6 74LS08
-23 -25 19 -17
0
0
13 VCC=14;GND=7;
0
0
0
5 DIP14
64

0 1 2 3 1 2 3 4 5 6
10 9 8 13 12 11 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0
0 0 0 0 4 1 2 0
1 U
7734 0 0
0
0
9 Inverter~
13 186 37 0 2 64
0 16 17
0
0 0 112 0
4 7404
-11 -20 17 -12
0
0
13 VCC=14;GND=7;
11 %D %1 %2 %S
0
0
5 DIP14
64

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0
88 0 0 0 6 1 1 0
1 U
9914 0 0
0
0
2 +V
167 55 143 0 1 64
0 3
0
0 0 53488 0
3 10V
-10 -22 11 -14
0
0
4 VCC;
10 %D %1 0 %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
7 Rocket~
180 569 302 0 20 64
20 4 2 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
-400
0
0 0 20528 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
9 Inverter~
13 366 218 0 2 64
0 8 5
0
0 0 112 0
4 7404
-11 -20 17 -12
0
0
13 VCC=14;GND=7;
11 %D %1 %2 %S
0
0
5 DIP14
64

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0
88 0 0 0 6 2 1 0
1 U
7931 0 0
0
0
12 SPST Switch~
165 488 312 0 2 64
0 4 5
0
0 0 20592 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
1 S
9325 0 0
0
0
13 Piezo Buzzer~
174 403 284 0 2 64
10 20 2
0
0 0 20528 270
0
0
0
0
0
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
12 2-Input AND~
0 372 250 0 3 64
0 8 21 20
0
0 0 48 0
6 74LS08
-23 -25 19 -17
0
0
13 VCC=14;GND=7;
0
0
0
5 DIP14
64

0 4 5 6 1 2 3 4 5 6
10 9 8 13 12 11 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0
0 0 0 0 4 2 2 0
1 U
3834 0 0
0
0
7 Ground~
168 403 338 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
8 Hex Key~
166 201 255 0 11 64
0 29 28 27 26 0 0 0 0 0
3 51
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -33686019
0 0 0 0 1 0 0 0
0
7668 0 0
0
0
6 74LS85
106 291 276 0 14 64
0 22 23 24 25 26 27 28 29 42
43 44 21 45 46
0
0 0 4272 0
6 74LS85
-21 -52 21 -44
0
0
13 VCC=16;GND=8;
0
0
0
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 -33686019
0 0 0 512 1 0 0 0
1 U
4718 0 0
0
0
7 Ground~
168 113 231 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3874 0 0
0
0
7 74LS168
8 159 154 0 30 64
0 2 2 19 3 2 2 3 16 2
8 22 23 24 25 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
9
0
0 0 4272 0
7 74LS168
-25 -61 24 -53
0
0
13 VCC=16;GND=8;
0
0
0
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 -33686019
0 0 0 0 1 0 0 0
1 U
6671 0 0
0
0
2 +V
167 406 17 0 1 64
0 3
0
0 0 53488 0
3 10V
-10 -22 11 -14
0
0
4 VCC;
10 %D %1 0 %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3789 0 0
0
0
9 CA 7-Seg~
184 406 71 0 18 64
10 15 14 13 12 11 10 9 2 3
0 0 0 2 2 0 0 0 1
0
0 0 20512 0
0
0
0
0
0
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 -33686019
0 0 0 0 1 0 0 0
0
4871 0 0
0
0
6 74LS47
187 288 147 0 14 64
0 22 23 24 25 47 48 9 10 11
12 13 14 15 49
0
0 0 4272 0
6 74LS47
-18 -61 24 -53
0
0
13 VCC=16;GND=8;
0
0
0
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 -33686019
0 0 0 512 1 0 0 0
1 U
3750 0 0
0
0
13 ResistorWire~
94 356 111 0 2 64
0 9 9
13 ResistorWire~
1 0 4112 0
0
0
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
0
8778 0 0
0
0
13 ResistorWire~
94 356 120 0 2 64
0 10 10
13 ResistorWire~
2 0 4112 0
0
0
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
0
538 0 0
0
0
13 ResistorWire~
94 356 129 0 2 64
0 11 11
13 ResistorWire~
3 0 4112 0
0
0
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
0
6843 0 0
0
0
13 ResistorWire~
94 356 138 0 2 64
0 12 12
13 ResistorWire~
4 0 4112 0
0
0
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
0
3136 0 0
0
0
13 ResistorWire~
94 356 147 0 2 64
0 13 13
13 ResistorWire~
5 0 4112 0
0
0
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
0
5950 0 0
0
0
13 ResistorWire~
94 356 156 0 2 64
0 14 14
13 ResistorWire~
6 0 4112 0
0
0
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
0
5670 0 0
0
0
13 ResistorWire~
94 356 165 0 2 64
0 15 15
13 ResistorWire~
7 0 4112 0
0
0
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
0
6828 0 0
0
0
9 Resistor~
219 15 185 0 4 64
0 6 3 0 1
9 Resistor~
0 0 4208 90
2 1k
-7 -28 7 -20
0
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
60
1 1 4 0 0 4224 0 9 11 0 0 2
537 312
505 312
2 2 5 0 0 8320 0 10 11 0 0 4
387 218
439 218
439 312
471 312
1 0 6 0 0 8320 0 2 0 0 15 4
39 118
5 118
5 210
15 210
3 1 7 0 0 12416 0 5 6 0 0 4
312 18
329 18
329 53
155 53
8 1 2 0 0 4096 0 20 1 0 0 2
427 107
427 125
2 0 3 0 0 8192 0 29 0 0 12 3
15 167
15 163
55 163
0 2 2 0 0 4096 0 0 2 14 0 2
113 118
73 118
0 4 8 0 0 4224 0 0 3 37 0 4
217 218
5 218
5 268
18 268
2 0 2 0 0 4224 0 9 0 0 10 2
537 321
403 321
2 1 2 0 0 0 0 12 14 0 0 2
403 315
403 332
4 0 3 0 0 4224 0 18 0 0 12 2
127 163
55 163
7 1 3 0 0 0 0 18 8 0 0 3
127 190
55 190
55 152
9 0 2 0 0 0 0 18 0 0 14 4
191 127
208 127
208 203
113 203
1 1 2 0 0 0 0 18 17 0 0 3
121 118
113 118
113 225
1 3 6 0 0 0 0 29 3 0 0 3
15 203
15 259
18 259
7 2 9 0 0 8320 0 20 22 0 0 3
421 107
421 111
374 111
2 6 10 0 0 4224 0 23 20 0 0 3
374 120
415 120
415 107
5 2 11 0 0 8320 0 20 24 0 0 3
409 107
409 129
374 129
2 4 12 0 0 8320 0 25 20 0 0 3
374 138
403 138
403 107
3 2 13 0 0 4224 0 20 26 0 0 3
397 107
397 147
374 147
2 2 14 0 0 8320 0 27 20 0 0 3
374 156
391 156
391 107
1 2 15 0 0 4224 0 20 28 0 0 3
385 107
385 165
374 165
1 13 15 0 0 0 0 28 21 0 0 2
338 165
326 165
12 1 14 0 0 0 0 21 27 0 0 2
326 156
338 156
1 11 13 0 0 0 0 26 21 0 0 2
338 147
326 147
10 1 12 0 0 0 0 21 25 0 0 2
326 138
338 138
1 9 11 0 0 0 0 24 21 0 0 2
338 129
326 129
8 1 10 0 0 0 0 21 23 0 0 2
326 120
338 120
1 7 9 0 0 0 0 22 21 0 0 2
338 111
326 111
1 0 16 0 0 8192 0 7 0 0 59 3
171 37
158 37
158 17
2 1 17 0 0 8320 0 7 4 0 0 4
207 37
217 37
217 72
209 72
0 2 8 0 0 0 0 0 4 37 0 3
217 154
217 84
209 84
3 2 18 0 0 8320 0 4 6 0 0 4
164 78
159 78
159 65
155 65
3 3 19 0 0 8320 0 6 18 0 0 4
110 59
103 59
103 136
127 136
3 1 20 0 0 4224 0 13 12 0 0 3
393 250
403 250
403 253
1 0 8 0 0 0 0 13 0 0 37 3
348 244
336 244
336 218
10 1 8 0 0 0 0 18 10 0 0 4
197 154
217 154
217 218
351 218
2 0 2 0 0 0 0 18 0 0 14 2
121 127
113 127
5 0 2 0 0 0 0 18 0 0 14 2
127 172
113 172
6 0 2 0 0 0 0 18 0 0 14 2
127 181
113 181
12 2 21 0 0 8320 0 16 13 0 0 4
323 294
335 294
335 256
348 256
1 4 22 0 0 4160 0 16 0 0 58 2
259 249
235 249
2 3 23 0 0 4160 0 16 0 0 58 2
259 258
235 258
3 2 24 0 0 4160 0 16 0 0 58 2
259 267
235 267
4 1 25 0 0 4160 0 16 0 0 58 2
259 276
235 276
5 4 26 0 0 4224 0 16 15 0 0 3
259 285
192 285
192 279
6 3 27 0 0 4224 0 16 15 0 0 3
259 294
198 294
198 279
7 2 28 0 0 4224 0 16 15 0 0 3
259 303
204 303
204 279
8 1 29 0 0 4224 0 16 15 0 0 3
259 312
210 312
210 279
4 1 25 0 0 0 0 21 0 0 58 2
256 138
235 138
3 2 24 0 0 0 0 21 0 0 58 2
256 129
235 129
2 3 23 0 0 0 0 21 0 0 58 2
256 120
235 120
4 1 22 0 0 0 0 0 21 58 0 2
235 111
256 111
14 1 25 0 0 4288 0 18 0 0 58 2
191 190
235 190
13 2 24 0 0 4288 0 18 0 0 58 2
191 181
235 181
12 3 23 0 0 4288 0 18 0 0 58 2
191 172
235 172
11 4 22 0 0 4288 0 18 0 0 58 2
191 163
235 163
2 0 1 0 0 4256 0 0 0 0 0 2
235 93
235 281
9 8 16 0 0 8320 0 3 18 0 0 6
88 250
94 250
94 17
225 17
225 118
197 118
1 9 3 0 0 0 0 19 20 0 0 2
406 26
406 35
4
-17 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 10
448 275 544 302
452 279 534 298
10 Arm/Safety
-17 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 21
434 48 537 98
438 52 527 90
21 Count down
to launch
-17 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 6
12 70 80 97
16 74 70 93
6 Launch
-17 0 0 0 700 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 14
109 252 188 302
113 256 178 294
14 Warning
Count
0
17 0 0
0
0
3 Vin
-1.5 -0.7 0.01
3 Vcc
10 14 1
100 0 1 100000
0 0.0005 2.5e-006 2.5e-006 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
0.00012 0.000100092 -7.7 -11.9 1.9908e-005 4.2
0 0
0 1 100
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
0.005 0 0.8 -0.4 0.005 0.005
16 0
0 0.001 100
0
0 0 100 100 0 0
98 66 294 126
0 0 0 0
294 66
98 66
294 66
294 126
0 0
19108.5 10 56 60.2 19098.5 19098.5
12387 0
0 5000 10000
0
0 0 100 100 0 0
77 66 293 126
0 0 0 0
293 66
77 66
293 66
293 126
0 0
1e+006 1 -3.55271e-015 -3.55271e-015 999999 999999
4211 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
