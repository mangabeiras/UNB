CircuitMaker Text
5.6
Probes: 2
charge
Transient Analysis
0 168 123 65280
discharge
Transient Analysis
1 386 117 65535
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
245 80 857 634
7 5.000 V
7 5.000 V
3 GND
2500 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
2 4 0.500000 0.500000
245 357 857 634
9961474 0
0
0
0
0
0
0
9
4 .IC~
207 366 89 0 1 64
0 3
0
0 0 53584 0
3 10v
-10 -16 11 -8
4 CMD1
-14 -26 14 -18
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
3 CMD
631 0 0
2
36626.4 0
0
7 Ground~
168 324 214 0 1 64
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
9466 0 0
2
36626.4 1
0
10 Capacitor~
219 397 154 0 2 64
0 2 3
10 Capacitor~
0 0 336 90
3 1uF
11 -5 32 3
2 C1
14 -15 28 -7
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
3266 0 0
2
36626.4 2
0
4 .IC~
207 149 93 0 1 64
0 4
0
0 0 53584 0
2 0V
-7 -16 7 -8
4 CMD2
-14 -26 14 -18
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
3 CMD
7693 0 0
2
36626.4 3
0
7 Ground~
168 107 218 0 1 64
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
3723 0 0
2
36626.4 4
0
10 Capacitor~
219 180 158 0 2 64
0 2 4
10 Capacitor~
0 0 336 90
3 1uF
11 -5 32 3
2 C2
14 -15 28 -7
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
3440 0 0
2
36626.4 5
0
8 Battery~
219 34 162 0 2 64
0 5 2
8 Battery~
0 0 368 0
3 10V
12 -7 33 1
2 V1
15 -17 29 -9
0
0
14 %D %1 %2 DC %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 -1 286 0 1 0 0 0
1 V
6263 0 0
2
36626.4 6
0
9 Resistor~
219 313 118 0 3 64
0 2 3 -1
9 Resistor~
0 0 368 0
3 200
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
4900 0 0
2
36626.4 7
0
9 Resistor~
219 96 122 0 2 64
0 5 4
9 Resistor~
0 0 368 0
3 200
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
8783 0 0
2
36626.4 8
0
9
1 0 3 0 0 4096 0 1 0 0 4 2
366 101
366 118
1 0 2 0 0 4096 0 2 0 0 3 2
324 208
324 190
1 1 2 0 0 8320 0 3 8 0 0 5
397 163
397 190
251 190
251 118
295 118
2 2 3 0 0 4224 0 8 3 0 0 3
331 118
397 118
397 145
1 0 4 0 0 4096 0 4 0 0 8 2
149 105
149 122
1 0 2 0 0 0 0 5 0 0 7 2
107 212
107 194
1 2 2 0 0 0 0 6 7 0 0 4
180 167
180 194
34 194
34 173
2 2 4 0 0 4224 0 9 6 0 0 3
114 122
180 122
180 149
1 1 5 0 0 8320 0 7 9 0 0 3
34 149
34 122
78 122
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 9
386 102 461 118
386 102 461 118
9 discharge
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 6
168 106 219 122
168 106 219 122
6 charge
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 172
8 4 504 68
12 8 500 56
172 Charging/Discharing capacitor example. The initial condition 
devices are required in order to make the capacitors start 
at the inital value of 0v or 10v respectively.
0
16 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.002 1.5e-05 1.5e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3952 8550464 100 100 0 0
77 66 977 276
0 403 1024 740
977 66
77 66
977 66
977 276
0 0
0 0 0 0 0 0
16 3
4 0.0005 5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
