CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 305 259
7 5.000 V
7 5.000 V
3 GND
2e+006 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 305 259
142606338 0
0
0
0
0
0
0
6
13 Logic Switch~
5 224 115 0 2 11
0 2 -99
0
0 0 4192 512
2 0V
-7 -16 7 -8
2 S1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 152 29 0 2 11
0 4 -99
0
0 0 4192 0
2 0V
-7 -16 7 -8
2 S2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 56 115 0 2 11
0 5 -99
0
0 0 4192 0
2 0V
-7 -16 7 -8
2 S3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 55 91 0 2 11
0 6 -99
0
0 0 4192 0
2 0V
-7 -16 7 -8
2 S4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
4 SIP3
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
4 LED~
171 177 65 0 2 5
10 4 3
0
0 0 96 0
4 LED2
10 -16 38 -8
2 D1
17 -26 31 -18
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5394 0 0
0
0
14 Opto Isolator~
173 136 103 0 4 9
0 6 5 3 2
0
0 0 96 0
6 OP4N25
-22 -28 20 -20
2 U1
-8 -38 6 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 -33686019
88 0 0 0 1 1 0 0
1 U
7734 0 0
0
0
5
1 4 2 0 0 4224 0 1 6 0 0 2
212 115
162 115
3 2 3 0 0 8320 0 6 5 0 0 3
162 91
177 91
177 75
1 1 4 0 0 8320 0 2 5 0 0 3
164 29
177 29
177 55
2 1 5 0 0 4224 0 6 3 0 0 2
108 115
68 115
1 1 6 0 0 4224 0 4 6 0 0 2
67 91
108 91
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 2.5e-006 1e-008 1e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3616 1210432 100 100 0 0
77 66 617 126
0 66 140 136
617 66
77 66
617 66
617 126
0 0
0 0 0 0 0 0
16 0
4 1 2
1
174 91
0 3 0 0 1	0 2 0 0
3412 8550464 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
0 0 0 0 0 0
0 0
4 5e-007 2
1
87 91
0 6 0 0 1	0 5 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
