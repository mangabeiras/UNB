CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 30 30 100 9
0 66 320 259
7 5.000 V
7 5.000 V
3 GND
16666.7 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 320 259
12058624 0
0
0
0
0
0
0
11
5 SAVE-
218 218 87 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
39 *Combine
*AC 0 1
*DC 7 12
*TRAN -1 1
0
0
0
1

0 0
0 0 0 0 1 0 0 0
4 SAVE
8953 0 0
0
0
5 SAVE-
218 97 109 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
20 *Combine
*TRAN -1 1
0
0
0
1

0 0
0 0 0 0 1 0 0 0
4 SAVE
4441 0 0
0
0
7 Ground~
168 218 176 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
2 +V
167 173 156 0 1 3
0 4
0
0 0 54112 180
4 -12V
-13 1 15 9
3 Vee
-10 11 11 19
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
2 +V
167 173 80 0 1 3
0 3
0
0 0 54112 0
4 +12V
-13 -14 15 -6
3 Vcc
-8 -24 13 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
7 Ground~
168 121 152 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
11 Signal Gen~
195 61 114 0 19 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 -1110651699 1176256512 0 1036831949
20
-0.1 10000 0 0.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -100m/100mV
-39 -30 38 -22
3 Vin
-11 -40 10 -32
0
0
44 %D %1 %2 DC 0 SIN(0 100m 10k 0 0) AC -100m 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
8 Op-Amp5~
219 173 115 0 5 11
0 2 5 3 4 6
8 Op-Amp5~
0 0 832 0
5 UA741
7 -15 42 -7
2 U1
17 -26 31 -18
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 -33686019
88 0 0 256 1 1 0 0
1 U
3747 0 0
0
0
9 Resistor~
219 218 143 0 3 5
0 2 6 -1
9 Resistor~
0 0 4960 90
3 25k
7 0 28 8
2 RL
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 185 50 0 2 5
0 5 6
9 Resistor~
0 0 4960 0
4 100k
-14 -12 14 -4
2 RF
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 121 109 0 2 5
0 7 5
9 Resistor~
0 0 4960 0
3 10k
-10 -12 11 -4
2 RI
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
9325 0 0
0
0
10
1 0 2 0 0 4096 0 6 0 0 2 2
121 146
121 121
1 2 2 0 0 4224 0 8 7 0 0 4
155 121
103 121
103 119
92 119
1 1 2 0 0 0 0 9 3 0 0 2
218 161
218 170
3 1 3 0 0 4224 0 8 5 0 0 2
173 102
173 89
4 1 4 0 0 4224 0 8 4 0 0 2
173 128
173 141
1 0 5 0 0 8320 0 10 0 0 7 3
167 50
147 50
147 109
2 2 5 0 0 0 0 11 8 0 0 2
139 109
155 109
2 0 6 0 0 8320 0 10 0 0 9 3
203 50
218 50
218 115
5 2 6 0 0 0 0 8 9 0 0 3
191 115
218 115
218 125
1 1 7 0 0 4224 0 7 11 0 0 2
92 109
103 109
0
0
29 0 1
0
0
3 Vin
-1.5 -0.7 0.02
3 Vcc
10 14 1
100 0 1 1e+006
0 0.0003 2.5e-006 2.5e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3588 1210432 100 100 0 0
98 66 608 126
0 66 140 136
608 66
77 66
617 66
617 126
0 0
5.34602e-315 1.57621e-314 5.18065e-315 1.56912e-314 5.34602e-315 5.18894e-315
0 0
4 1 5
1
173 95
0 3 0 0 1	0 4 0 0
3684 8550976 100 100 0 0
77 66 287 126
0 259 320 452
287 66
77 66
287 66
287 126
0 0
4.77568e-315 0 5.27183e-315 1.58818e-314 4.77568e-315 4.77568e-315
121 0
4 0.0001 5
1
218 81
0 6 0 0 2	0 8 0 0
4052 2259008 100 100 0 0
77 66 287 126
320 66 640 259
287 66
77 66
287 66
287 126
0 0
1.58503e-314 1.58942e-314 5.41171e-315 5.37959e-315 5.24531e-315 5.24531e-315
0 0
4 0.3 1e+036
1
218 74
0 6 0 0 2	0 8 0 0
3700 4421696 100 100 0 0
77 66 293 126
320 259 640 452
293 66
77 66
293 66
293 66
0 0
6.08861e-315 5.26354e-315 1.38842e-314 1.38842e-314 6.08861e-315 6.08861e-315
4211 0
4 300000 500000
1
218 78
0 6 0 0 2	0 8 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
