CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 36 30 100 3
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
0 66 640 259
9961474 0
0
0
0
0
0
0
14
7 Trans2~
219 159 115 0 4 9
0 8 2 7 6
0
0 0 336 0
5 10TO1
-16 -32 19 -24
2 T1
-6 -42 8 -34
0
0
17 %D %1 %2 %3 %4 %S
0
24 alias:XTRANS {RATIO=0.1}
0
9

0 1 2 3 4 1 2 3 4 0
88 0 0 0 1 0 0 0
1 T
8953 0 0
0
0
5 SAVE-
218 490 75 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
20 *Combine
*TRAN 0 16
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SAVE-
218 310 75 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
20 *Combine
*TRAN 0 16
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SAVE-
218 113 104 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 C
3 -26 10 -18
0
0
0
14 *TRAN -170 170
0
0
0
1

0 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
7 Ground~
168 561 186 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 106 158 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
11 Signal Gen~
195 49 114 0 19 64
0 8 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1114636288 0 1126825984
20
1 60 0 170 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 17232 0
9 -170/170V
-31 -28 32 -20
2 V1
-7 -38 7 -30
0
0
38 %D %1 %2 DC 0 SIN(0 170 60 0 0) AC 1 0
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
10 FW Bridge~
219 252 123 0 4 9
0 2 7 5 6
10 FW Bridge~
0 0 848 0
6 18DB10
-17 -57 25 -49
2 D1
-4 -67 10 -59
0
0
17 %D %1 %2 %3 %4 %S
0
0
3 D-2
9

0 1 2 3 4 1 2 3 4 0
88 0 0 256 1 0 0 0
1 D
3747 0 0
0
0
10 Polar Cap~
219 330 122 0 2 5
0 5 2
10 Polar Cap~
0 0 848 270
5 100uF
10 4 45 12
2 C1
21 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
3549 0 0
0
0
12 Zener Diode~
219 437 149 0 2 5
0 2 4
12 Zener Diode~
0 0 848 90
6 1N4736
14 -2 56 6
2 D2
28 -12 42 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
100 0 0 0 1 1 0 0
1 D
7931 0 0
0
0
12 NPN Trans:C~
219 441 82 0 3 7
0 5 4 3
12 NPN Trans:C~
0 0 848 90
7 2N2222A
-27 -26 22 -18
2 Q1
-9 -36 5 -28
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 -33686019
81 0 0 0 1 1 0 0
1 Q
9325 0 0
0
0
10 Polar Cap~
219 505 123 0 2 5
0 3 2
10 Polar Cap~
0 0 848 26894
5 100uF
10 4 45 12
2 C2
21 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
8903 0 0
0
0
9 Resistor~
219 389 101 0 2 64
0 5 4
9 Resistor~
0 0 4976 270
3 680
7 1 28 9
2 R1
8 -11 22 -3
0
0
11 %D %1 %2 %V
0
0
0
3

0 1 2 1
82 0 0 0 1 1 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 561 115 0 3 5
0 2 3 -1
9 Resistor~
0 0 4976 90
2 5k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3363 0 0
0
0
17
2 0 2 0 0 4096 0 12 0 0 16 2
504 130
504 169
1 0 3 0 0 4096 0 12 0 0 6 2
504 113
504 75
2 0 4 0 0 8320 0 13 0 0 5 3
389 119
389 126
439 126
1 0 5 0 0 4096 0 13 0 0 17 2
389 83
389 75
2 2 4 0 0 0 0 11 10 0 0 2
439 98
439 137
3 2 3 0 0 4224 0 11 14 0 0 3
457 75
561 75
561 97
1 0 2 0 0 0 0 6 0 0 10 2
106 152
106 126
4 4 6 0 0 8320 0 8 1 0 0 5
254 151
254 159
185 159
185 134
177 134
3 2 7 0 0 12416 0 1 8 0 0 5
177 96
187 96
187 77
254 77
254 87
2 2 2 0 0 4096 0 1 7 0 0 3
141 126
80 126
80 119
1 1 8 0 0 4224 0 1 7 0 0 3
141 104
80 104
80 109
2 0 2 0 0 0 0 9 0 0 16 2
329 129
329 169
1 0 5 0 0 4096 0 9 0 0 17 2
329 112
329 75
1 0 2 0 0 0 0 14 0 0 16 2
561 133
561 169
1 0 2 0 0 0 0 10 0 0 16 2
439 157
439 169
1 1 2 0 0 12416 0 8 5 0 0 5
222 119
215 119
215 169
561 169
561 180
3 1 5 0 0 12416 0 8 11 0 0 4
286 119
295 119
295 75
421 75
1
-16 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 20
217 5 427 34
222 9 422 28
20 +6 Volt Power Supply
35 .OPTIONS ABSTOL=1.000u ITL4=100.0

16 0 0
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 0.08333 0.0004167 0.0004167 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
2140 8550976 100 100 0 0
98 66 608 126
0 259 640 452
608 66
98 66
608 71
608 116
0 0
0.08333 0 18 0 0.08333 0.08333
12409 0
4 0.02 100
3
339 75
0 5 0 0 3	0 17 0 0
213 77
0 7 0 0 3	0 9 0 0
493 75
0 3 0 0 1	0 6 0 0
0 0 100 100 0 0
77 66 617 126
0 0 0 0
617 66
77 66
617 66
617 126
0 0
0.0003 0 5 0 0.0003 0.0003
13433 0
0 5e-005 5
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
-0.72 -1.5 12.6 7.2 0.78 0.78
0 0
0 0.3 1e+036
0
0 0 100 100 0 0
77 66 293 126
0 0 0 0
293 66
77 66
293 66
293 126
0 0
1e+006 1 -3.55271e-015 -3.55271e-015 999999 999999
4211 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
