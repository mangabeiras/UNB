CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 18 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
0 66 320 452
7 5.000 V
7 5.000 V
3 GND
41666.7 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 320 452
12058632 0
0
0
0
0
0
0
18
5 SAVE-
218 343 150 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
31 *Combine
*AC -1 25
*TRAN -5 5
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 78 183 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
20 *Combine
*TRAN -5 5
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
7 Ground~
168 357 215 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
7 Ground~
168 215 283 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
7 Ground~
168 73 219 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
11 Signal Gen~
195 32 188 0 19 64
0 9 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1036831949 1209810944 0 1008981770
20
0.1 160000 0 0.01 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
9 -10m/10mV
-31 -28 32 -20
2 V1
-7 -38 7 -30
0
0
43 %D %1 %2 DC 0 SIN(0 10m 160k 0 0) AC 100m 0
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
2 +V
167 215 24 0 1 64
0 7
0
0 0 54112 0
4 -10V
13 -4 41 4
3 Vcc
-9 -17 12 -9
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
12 PNP Trans:C~
219 210 183 0 3 64
0 3 5 8
12 PNP Trans:C~
0 0 320 0
6 2N3906
20 -4 62 4
2 Q1
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
113 0 0 0 1 0 0 0
1 Q
3747 0 0
0
0
8 Coil 3T~
219 215 74 0 2 64
0 6 7
8 Coil 3T~
0 0 832 90
4 96uH
8 -4 36 4
2 LT
9 -15 23 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
76 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
10 Capacitor~
219 265 97 0 2 64
0 3 7
10 Capacitor~
0 0 832 90
5 .01uF
9 2 44 10
2 CT
15 -9 29 -1
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
7931 0 0
0
0
10 Capacitor~
219 265 239 0 2 64
0 2 8
10 Capacitor~
0 0 832 90
4 15uF
14 2 42 10
2 CE
14 -9 28 -1
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
9325 0 0
0
0
10 Capacitor~
219 105 183 0 2 64
0 9 5
10 Capacitor~
0 0 832 0
5 .03uF
-14 -20 21 -12
2 Ci
-5 -31 9 -23
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
8903 0 0
0
0
10 Capacitor~
219 313 150 0 2 64
0 3 4
10 Capacitor~
0 0 832 0
5 .03uF
-18 -18 17 -10
2 Co
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3834 0 0
0
0
9 Resistor~
219 133 104 0 4 64
0 5 7 0 1
9 Resistor~
0 0 864 90
3 18k
8 0 29 8
2 R1
11 -11 25 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 133 241 0 3 64
0 2 5 -1
9 Resistor~
0 0 864 90
3 33k
7 2 28 10
2 R2
8 -9 22 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 215 238 0 3 64
0 2 8 -1
9 Resistor~
0 0 864 90
2 1k
7 2 21 10
2 RE
7 -9 21 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 215 121 0 2 64
0 3 6
9 Resistor~
0 0 864 90
3 6.3
8 -1 29 7
2 Rs
8 -12 22 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 357 179 0 3 64
0 2 4 -1
9 Resistor~
0 0 864 90
3 10k
8 1 29 9
2 RL
10 -10 24 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
19
1 0 3 0 0 4096 0 13 0 0 7 2
304 150
265 150
2 2 4 0 0 4224 0 13 18 0 0 3
322 150
357 150
357 161
1 1 2 0 0 4096 0 18 3 0 0 2
357 197
357 209
1 0 5 0 0 4096 0 14 0 0 6 2
133 122
133 183
2 0 5 0 0 0 0 15 0 0 6 2
133 223
133 183
2 2 5 0 0 4224 0 12 8 0 0 2
114 183
192 183
1 0 3 0 0 8320 0 10 0 0 8 3
265 106
265 150
215 150
1 1 3 0 0 0 0 17 8 0 0 2
215 139
215 165
1 2 6 0 0 4224 0 9 17 0 0 2
215 94
215 103
2 0 7 0 0 8320 0 14 0 0 14 3
133 86
133 42
215 42
2 0 7 0 0 0 0 10 0 0 14 3
265 88
265 42
215 42
1 0 2 0 0 8192 0 11 0 0 18 3
265 248
265 268
215 268
2 0 8 0 0 8320 0 11 0 0 17 3
265 230
265 212
215 212
1 2 7 0 0 0 0 7 9 0 0 2
215 33
215 54
2 1 2 0 0 0 0 6 5 0 0 3
63 193
73 193
73 213
1 0 2 0 0 0 0 4 0 0 18 2
215 277
215 268
2 3 8 0 0 0 0 16 8 0 0 2
215 220
215 201
1 1 2 0 0 8320 0 15 16 0 0 4
133 259
133 268
215 268
215 256
1 1 9 0 0 4224 0 6 12 0 0 2
63 183
96 183
1
-16 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 18
5 9 195 38
9 13 189 32
18 Bandpass Amplifier
0
24 0 1
0
0
0
0 0 0
0
0 0 0
200 1 10000 1e+006
0.0001 0.00012 1.5e-007 1.5e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3496 8550464 100 100 0 0
77 66 287 126
320 66 640 259
287 66
77 66
287 66
287 126
0 0
4.72335e-315 4.70983e-315 1.59948e-314 1.60181e-314 4.61305e-315 4.61305e-315
16 0
4 3e-005 5
1
281 150
0 3 0 0 1	0 1 0 0
1948 4356160 100 100 0 0
77 66 297 126
320 259 640 452
297 66
77 66
297 66
297 126
0 0
6.08861e-315 5.81148e-315 5.45005e-315 0 6.08782e-315 6.08782e-315
18 0
4 300000 500000
1
284 150
0 3 0 0 1	0 1 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
