CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
16 4 30 100 3
16 82 362 310
7 5.000 V
7 5.000 V
3 GND
16 82 362 310
9437184 0
0
0
0
0
0
0
6
13 Logic Switch~
5 183 116 0 2 3
0 2 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
0
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
8 Hex Key~
166 125 58 0 11 11
0 3 4 5 6 0 0 0 0 0
0 48
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4441 0 0
0
0
12 Hex Display~
7 292 62 0 4 9
10 3 4 5 6
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
0
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3618 0 0
0
0
14 Logic Display~
6 39 78 0 1 3
10 2
0
0 0 53344 0
6 100MEG
3 -16 45 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
11 DB-9 Macro~
94 242 134 0 9 19
0 10 9 8 7 2 3 4 5 6
11 DB-9 Macro~
1 0 4112 0
0
0
0
0
0
0
0
0
19

0 0 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451
0 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
11 DB-9 Macro~
94 80 134 0 9 19
0 10 9 8 7 2 3 4 5 6
11 DB-9 Macro~
2 0 4112 0
0
0
0
0
0
0
0
0
19

0 0 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451
0 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451 -842150451 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
10
1 5 2 0 0 4224 0 1 5 0 0 2
195 116
220 116
1 5 2 0 0 0 0 4 6 0 0 3
39 96
39 116
58 116
6 1 3 0 0 8192 0 5 3 0 0 3
264 147
301 147
301 86
2 7 4 0 0 4096 0 3 5 0 0 3
295 86
295 138
264 138
8 3 5 0 0 8192 0 5 3 0 0 3
264 129
289 129
289 86
4 9 6 0 0 4096 0 3 5 0 0 3
283 86
283 120
264 120
1 6 3 0 0 4224 0 2 6 0 0 3
134 82
134 147
102 147
2 7 4 0 0 4224 0 2 6 0 0 3
128 82
128 138
102 138
3 8 5 0 0 4224 0 2 6 0 0 3
122 82
122 129
102 129
4 9 6 0 0 4224 0 2 6 0 0 3
116 82
116 120
102 120
0
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
0.002 0 0.09 -0.09 0.002 0.002
16 0
0 0.0005 10
0
0 0 100 100 0 0
98 66 294 126
0 0 0 0
294 66
98 66
294 66
294 126
0 0
1e+007 1 12.16 12.184 1e+007 1e+007
12403 0
0 3e+006 5e+006
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
2000 1 2.38857 0 1999 1999
16 0
0 500 1000
0
0 0 100 100 0 0
98 66 296 126
0 0 0 0
296 66
98 66
296 66
296 126
0 0
1e+006 1 -3.55271e-015 0 999999 999999
12403 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
