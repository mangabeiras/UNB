CircuitMaker Text
5.6
Probes: 15
U5_4
AC Analysis
2 466 136 16776960
U5_4
DC Sweep
2 466 136 16776960
U5_4
Operating Point
2 466 136 16776960
U5_4
Fourier Analysis
2 466 136 16776960
U5_5
AC Analysis
1 464 101 65535
U5_5
DC Sweep
1 464 101 65535
U5_5
Operating Point
1 464 101 65535
U5_5
Fourier Analysis
1 464 101 65535
U5_6
AC Analysis
0 439 92 65280
U5_6
DC Sweep
0 439 92 65280
U5_6
Operating Point
0 439 92 65280
U5_6
Fourier Analysis
0 439 92 65280
Q1
Transient Analysis
0 464 135 65280
Q2
Transient Analysis
1 464 100 65535
Q3
Transient Analysis
2 464 65 16776960
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 16 20 
10 13 13 10 20 13 46 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 15 100 10
231 152 911 669
8  5.000 V
8  5.000 V
3 GND
333333 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
2 4 0.386847 0.500000
231 469 911 669
11010050 0
0
0
0
0
0
0
21
7 Ground~
168 471 37 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8921 0 0
2
36626.6 3
0
7 74LS173
129 395 83 0 14 29
0 2 2 2 6 11 10 9 2 2
2 5 4 3 8
0
0 0 12528 0
7 74LS173
-24 -51 25 -43
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 -33686019
65 0 0 0 1 1 0 0
1 U
5910 0 0
2
36626.6 4
0
7 Ground~
168 427 230 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7815 0 0
2
36626.6 5
0
7 Ground~
168 592 149 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8481 0 0
2
36626.6 6
0
2 +V
167 592 35 0 1 3
0 12
0
0 0 53744 0
2 5V
-7 -22 7 -14
2 V1
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6241 0 0
2
36626.6 7
0
7 Ground~
168 279 81 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3972 0 0
2
36626.6 8
0
11 Signal Gen~
195 218 60 0 64 64
0 6 2 1 86 -9 9 0 0 0
0 0 0 0 0 0 0 1232348160 0 1084227584
869711765 841731191 841731191 869711765 897988541 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
20
0 1e+06 0 5 1e-07 1e-08 1e-08 1e-07 1e-06 0
0 0 0 0 0 0 0 0 0 0
0
0 0 16720 0
4 0/5V
-14 -28 14 -20
2 V2
-7 -38 7 -30
0
0
45 %D %1 %2 DC 0 PULSE(0 5 100n 10n 10n 100n 1u)
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
551 0 0
2
36626.6 9
0
9 Inverter~
13 518 136 0 2 21
0 3 13
0
0 0 368 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 1 1 0
1 U
4680 0 0
2
36626.6 10
0
9 Inverter~
13 518 101 0 2 21
0 4 7
0
0 0 368 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 2 1 0
1 U
8751 0 0
2
36626.6 11
0
9 Inverter~
13 518 65 0 2 21
0 5 11
0
0 0 368 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 3 1 0
1 U
9317 0 0
2
36626.6 12
0
8 2-In OR~
219 305 169 0 3 21
0 14 18 9
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 U2A
-2 -25 19 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 2 0
1 U
3481 0 0
2
36626.6 13
0
8 2-In OR~
219 237 160 0 3 21
0 16 15 14
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 U2B
-3 -24 18 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 2 2 0
1 U
6213 0 0
2
36626.6 14
0
8 2-In OR~
219 240 101 0 3 21
0 20 19 10
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 U2C
3 -24 24 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 3 2 0
1 U
3226 0 0
2
36626.6 15
0
9 2-In AND~
219 116 237 0 3 21
0 11 3 17
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U4C
-14 -25 7 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 3 6 0
1 U
7407 0 0
2
36626.6 16
0
9 2-In AND~
219 117 192 0 3 21
0 4 5 15
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U4B
-15 -24 6 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 2 6 0
1 U
9465 0 0
2
36626.6 17
0
9 2-In AND~
219 116 151 0 3 21
0 4 13 16
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -23 9 -15
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 6 0
1 U
4581 0 0
2
36626.6 18
0
9 2-In AND~
219 117 110 0 3 21
0 5 3 19
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U3B
-14 -24 7 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 2 5 0
1 U
3204 0 0
2
36626.6 19
0
9 2-In AND~
219 116 68 0 3 21
0 11 13 20
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U3A
-14 -24 7 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 1 5 0
1 U
9635 0 0
2
36626.6 20
0
9 2-In AND~
219 254 246 0 3 21
0 17 7 18
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U4D
-15 -25 6 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 -33686019
65 0 0 0 4 4 6 0
1 U
4377 0 0
2
36626.6 21
0
9 Resistor~
219 427 190 0 4 5
0 8 2 0 -1
0
0 0 368 270
3 10k
-30 -2 -9 6
2 R1
-27 -11 -13 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3672 0 0
2
36626.6 22
0
9 Resistor~
219 592 93 0 2 5
0 12 2
0
0 0 368 270
2 1k
8 -5 22 3
2 R2
7 -16 21 -8
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
8807 0 0
2
36626.6 23
0
36
8 0 2 0 0 8192 0 2 0 0 15 4
363 119
357 119
357 217
427 217
1 0 2 0 0 0 0 2 0 0 6 2
363 56
339 56
10 0 2 0 0 0 0 2 0 0 6 3
433 65
443 65
443 31
9 0 2 0 0 0 0 2 0 0 6 2
433 56
433 31
2 0 2 0 0 0 0 2 0 0 6 2
357 65
339 65
1 3 2 0 0 4224 0 1 2 0 0 4
471 31
339 31
339 74
357 74
1 4 6 0 0 4224 0 7 2 0 0 4
249 55
307 55
307 83
363 83
2 1 2 0 0 0 0 7 6 0 0 3
249 65
279 65
279 75
2 2 7 0 0 12416 0 9 19 0 0 6
539 101
556 101
556 268
217 268
217 255
230 255
11 1 5 0 0 12288 0 2 10 0 0 4
427 92
455 92
455 65
503 65
14 1 8 0 0 4224 0 2 20 0 0 2
427 119
427 172
7 3 9 0 0 8320 0 2 11 0 0 4
363 110
348 110
348 169
338 169
6 3 10 0 0 4224 0 2 13 0 0 2
363 101
273 101
5 0 11 0 0 8192 0 2 0 0 20 3
363 92
322 92
322 10
1 2 2 0 0 0 0 3 20 0 0 2
427 224
427 208
2 1 2 0 0 0 0 21 4 0 0 2
592 111
592 143
1 1 12 0 0 4224 0 5 21 0 0 2
592 44
592 75
2 2 13 0 0 12432 0 8 18 0 0 6
539 136
545 136
545 276
35 276
35 77
92 77
1 12 4 0 0 4096 0 9 2 0 0 2
503 101
427 101
2 1 11 0 0 12416 0 10 14 0 0 6
539 65
555 65
555 10
10 10
10 228
92 228
1 3 14 0 0 4224 0 11 12 0 0 2
292 160
270 160
2 3 15 0 0 4224 0 12 15 0 0 4
224 169
178 169
178 192
138 192
1 3 16 0 0 4224 0 12 16 0 0 2
224 151
137 151
1 3 17 0 0 4224 0 19 14 0 0 2
230 237
137 237
3 2 18 0 0 8320 0 19 11 0 0 4
275 246
281 246
281 178
292 178
2 0 3 0 0 4096 0 14 0 0 30 2
92 246
59 246
2 0 5 0 0 12416 0 15 0 0 10 5
93 201
22 201
22 18
455 18
455 65
1 0 4 0 0 0 0 15 0 0 35 2
93 183
70 183
2 0 13 0 0 0 0 16 0 0 18 2
92 160
35 160
2 13 3 0 0 12416 0 17 2 0 0 6
93 119
59 119
59 286
442 286
442 110
427 110
1 0 5 0 0 0 0 17 0 0 27 2
93 101
22 101
1 0 11 0 0 0 0 18 0 0 20 2
92 59
10 59
3 2 19 0 0 4224 0 17 13 0 0 2
138 110
227 110
3 1 20 0 0 12416 0 18 13 0 0 4
137 68
179 68
179 92
227 92
0 1 4 0 0 8320 0 0 16 19 0 5
455 101
455 296
70 296
70 142
92 142
0 1 3 0 0 0 0 0 8 30 0 2
442 136
503 136
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
469 120 488 136
469 120 488 136
2 Q1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
468 85 487 101
468 85 487 101
2 Q2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
467 49 486 65
467 49 486 65
2 Q3
44 .OPTIONS METHOD=GEAR MAXORD=2 GMINSTEP=100

16 0 0
0
0
3 Vin
-0.1 0.1 0.005
3 Vee
-15 0 1
100 0 1 1e+06
0 1.5e-05 1e-07 5e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
4016 8550976 100 100 0 0
77 66 617 276
0 417 652 768
617 66
77 66
617 66
617 276
0 0
0 0 0 0 0 0
5177 0
2 3e-06 3
3
442 120
10 18 0 -99 4	0 30 0 0
466 101
14 12 0 -21 1	0 19 0 0
455 82
16 5 0 47 2	0 10 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
