CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 15 100 9
0 66 530 437
7 5.000 V
7 5.000 V
3 GND
156250 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 530 437
143654914 0
0
0
0
0
0
0
12
9 Data Seq~
170 86 274 0 17 21
0 21 22 23 24 25 26 27 5 28
29 7 1 32 3 2 0 33
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -54 10 -46
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 DIP14
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
8953 0 0
0
0
AAAAABAAABAAABAAABAAABAAABAAABAAABAAABAAABAAABAAABAAABAAABAAABAAAB
7 Ground~
168 183 220 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
6 74LS75
103 101 108 0 14 29
0 9 10 5 11 4 5 3 30 6
31 7 32 8 33
0
0 0 12512 0
6 74LS75
-21 -51 21 -43
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
113 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 6 4 3 2 13 9 8 10
11 15 14 16 1 7 6 4 3 2
13 9 8 10 11 15 14 16 1 -33686019
65 0 0 512 1 1 0 0
1 U
3618 0 0
0
0
6 74LS93
109 105 197 0 8 17
0 2 2 5 4 9 10 11 4
0
0 0 12512 512
6 74LS93
-21 -35 21 -27
2 U2
-7 -45 7 -37
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 -33686019
65 0 0 0 1 1 0 0
1 U
6153 0 0
0
0
6 PROM32
80 201 108 0 14 29
0 2 2 3 6 7 8 34 35 36
37 15 14 13 12
0
0 0 12512 0
6 PROM32
-21 -19 21 -11
2 U3
-7 -29 7 -21
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 -33686019
65 0 0 512 1 1 0 0
1 U
5394 0 0
0
0
AKALAJANAFAHAGAOAKAOAGAHAFANAJALAKAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
8 Stepper~
185 422 92 0 6 13
13 20 16 19 18 16 17
0
0 0 4192 0
4 100H
10 -16 38 -8
2 M1
17 -26 31 -18
0
0
130 %DA %1 N%DA %V
R%DA N%DA %2 10
%DB %3 N%DB %V
R%DB N%DB %2 10
%DC %4 N%DC %V
R%DC N%DC %5 10
%DD %6 N%DD %V
R%DD N%DD %5 10
0
0
4 SIP6
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
76 0 0 0 1 0 0 0
1 M
7734 0 0
0
0
2 +V
167 486 60 0 1 3
0 16
0
0 0 53472 0
3 10V
12 -2 33 6
2 B1
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
7 Ground~
168 355 276 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
14 Opto Isolator~
173 316 217 0 10 64
0 12 2 17 2 0 0 0 0 0
10
0
0 0 96 0
7 OPTOISO
-26 -28 23 -20
2 U4
-9 -38 5 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
5

0 1 2 3 4 0
88 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
14 Opto Isolator~
173 316 169 0 10 64
0 13 2 18 2 0 0 0 0 0
10
0
0 0 96 0
7 OPTOISO
-26 -28 23 -20
2 U5
-9 -38 5 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
5

0 1 2 3 4 0
88 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
14 Opto Isolator~
173 316 120 0 10 64
0 14 2 19 2 0 0 0 0 0
10
0
0 0 96 0
7 OPTOISO
-26 -28 23 -20
2 U6
-9 -38 5 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
5

0 1 2 3 4 0
88 0 0 0 1 0 0 0
1 U
9325 0 0
0
0
14 Opto Isolator~
173 315 74 0 10 64
0 15 2 20 2 0 0 0 0 0
10
0
0 0 96 0
7 OPTOISO
-26 -28 23 -20
2 U7
-9 -38 5 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
5

0 1 2 3 4 0
88 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
34
2 0 2 0 0 4096 0 5 0 0 2 2
169 108
153 108
1 0 2 0 0 8192 0 5 0 0 5 3
163 72
153 72
153 188
7 3 3 0 0 8320 0 3 5 0 0 4
133 81
163 81
163 117
169 117
0 4 4 0 0 8320 0 0 4 15 0 5
46 215
46 231
146 231
146 215
137 215
2 0 2 0 0 0 0 4 0 0 6 3
131 197
153 197
153 188
1 1 2 0 0 0 0 4 2 0 0 3
131 188
183 188
183 214
6 0 5 0 0 4096 0 3 0 0 8 2
69 135
55 135
3 0 5 0 0 12416 0 3 0 0 16 5
69 99
55 99
55 165
161 165
161 206
4 9 6 0 0 8320 0 5 3 0 0 4
169 126
159 126
159 99
133 99
11 5 7 0 0 12416 0 3 5 0 0 4
133 117
147 117
147 135
169 135
13 6 8 0 0 12416 0 3 5 0 0 4
133 135
143 135
143 144
169 144
5 1 9 0 0 8320 0 4 3 0 0 4
67 188
14 188
14 81
69 81
2 6 10 0 0 8320 0 3 4 0 0 4
69 90
24 90
24 197
67 197
7 4 11 0 0 8320 0 4 3 0 0 4
67 206
35 206
35 117
69 117
5 8 4 0 0 0 0 3 4 0 0 4
69 126
46 126
46 215
67 215
8 3 5 0 0 0 0 1 4 0 0 4
118 310
161 310
161 206
137 206
14 1 12 0 0 8320 0 5 9 0 0 4
233 144
248 144
248 205
288 205
13 1 13 0 0 12416 0 5 10 0 0 4
233 135
254 135
254 157
288 157
12 1 14 0 0 12416 0 5 11 0 0 4
233 126
254 126
254 108
288 108
11 1 15 0 0 8320 0 5 12 0 0 4
233 117
248 117
248 62
287 62
1 0 16 0 0 4096 0 7 0 0 22 3
486 69
486 92
465 92
2 5 16 0 0 8320 0 6 6 0 0 4
458 68
465 68
465 116
458 116
2 0 2 0 0 0 0 11 0 0 26 2
288 132
262 132
2 0 2 0 0 0 0 10 0 0 26 2
288 181
262 181
2 0 2 0 0 0 0 9 0 0 26 2
288 229
262 229
2 0 2 0 0 8192 0 12 0 0 34 4
287 86
262 86
262 254
355 254
3 6 17 0 0 8320 0 9 6 0 0 4
342 205
379 205
379 122
386 122
3 4 18 0 0 8320 0 10 6 0 0 4
342 157
372 157
372 110
386 110
3 3 19 0 0 8320 0 11 6 0 0 4
342 108
365 108
365 74
386 74
3 1 20 0 0 4224 0 12 6 0 0 2
341 62
386 62
4 0 2 0 0 0 0 11 0 0 34 2
342 132
355 132
4 0 2 0 0 0 0 10 0 0 34 2
342 181
355 181
4 0 2 0 0 0 0 9 0 0 34 2
342 229
355 229
4 1 2 0 0 8320 0 12 8 0 0 3
341 86
355 86
355 270
4
-13 0 0 0 700 0 0 0 0 3 2 1 34
5 Arial
0 0 0 14
391 1 448 42
395 5 445 37
14 Stepper
Motor
-13 0 0 0 700 0 0 0 0 3 2 1 34
5 Arial
0 0 0 16
284 3 354 44
288 7 351 39
16 Opto-
Isolators
-13 0 0 0 700 0 0 0 0 3 2 1 34
5 Arial
0 0 0 4
176 4 222 26
180 8 219 24
4 PROM
-13 0 0 0 700 0 0 0 0 3 2 1 34
5 Arial
0 0 0 20
68 3 142 44
72 7 139 39
20 Counter & 
Latches
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 3.2e-005 1.28e-007 1.28e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3224 8525888 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
0 0 0 0 0 0
16 0
4 1e-005 100
1
360 62
0 20 0 0 1	0 30 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
