CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 100 9
0 66 640 259
8  5.000 V
8  5.000 V
3 GND
5000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 259
9961488 0
0
0
0
0
0
0
11
5 SAVE-
218 38 115 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
11 *TRAN -1 13
0
3 0�t
0
1

0 0
0 0 0 0 1 0 0 0
4 SAVE
8953 0 0
0
0
4 .IC~
207 98 144 0 1 3
0 4
0
0 0 53312 0
2 0V
-7 -15 7 -7
2 V2
-7 -25 7 -17
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
3 CMD
4441 0 0
0
0
2 +V
167 166 37 0 1 3
0 6
0
0 0 53600 0
4 +12V
9 -2 37 6
2 V1
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
10 555 Timer~
219 108 106 0 8 17
0 2 4 8 7 5 4 3 6
10 555 Timer~
0 0 6464 0
3 555
-10 -23 11 -15
2 U1
-7 -33 7 -25
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 -33686019
88 0 0 0 1 1 0 0
1 U
6153 0 0
0
0
10 Polar Cap~
219 213 187 0 2 5
0 4 2
10 Polar Cap~
0 0 832 26894
4 .1uF
8 4 36 12
2 CT
16 -6 30 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
5394 0 0
0
0
10 Polar Cap~
219 160 186 0 2 5
0 5 2
10 Polar Cap~
0 0 832 26894
5 .01uF
5 4 40 12
2 C1
21 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
7734 0 0
0
0
7 Ground~
168 112 227 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
9 Resistor~
219 14 157 0 3 5
0 2 8 -1
9 Resistor~
0 0 4960 90
3 10k
7 0 28 8
2 RL
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 212 73 0 4 5
0 3 6 0 1
9 Resistor~
0 0 4960 90
2 1k
8 0 22 8
2 RA
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 212 133 0 2 5
0 4 3
9 Resistor~
0 0 4960 90
2 1k
8 0 22 8
2 RB
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 29 81 0 4 5
0 7 6 0 1
9 Resistor~
0 0 4960 90
2 2k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
9325 0 0
0
0
16
2 0 3 0 0 4096 0 10 0 0 2 2
212 115
212 106
7 1 3 0 0 4224 0 4 9 0 0 3
140 106
212 106
212 91
1 0 4 0 0 4096 0 2 0 0 13 2
98 156
98 164
2 0 2 0 0 4096 0 6 0 0 11 2
159 193
159 206
1 5 5 0 0 4224 0 6 4 0 0 3
159 176
159 124
140 124
1 0 2 0 0 4096 0 7 0 0 11 2
112 221
112 206
2 0 6 0 0 8320 0 11 0 0 16 3
29 63
29 60
166 60
4 1 7 0 0 4224 0 4 11 0 0 3
76 124
29 124
29 99
1 0 2 0 0 8192 0 8 0 0 11 3
14 175
14 186
51 186
3 2 8 0 0 4224 0 4 8 0 0 3
76 115
14 115
14 139
1 2 2 0 0 12416 0 4 5 0 0 5
76 97
51 97
51 206
212 206
212 194
1 0 4 0 0 4096 0 5 0 0 14 2
212 177
212 164
2 0 4 0 0 12416 0 4 0 0 14 4
76 106
65 106
65 164
185 164
6 1 4 0 0 0 0 4 10 0 0 5
140 115
185 115
185 164
212 164
212 151
2 0 6 0 0 0 0 9 0 0 16 3
212 55
212 51
166 51
1 8 6 0 0 0 0 3 4 0 0 3
166 46
166 97
140 97
0
27 .OPTIONS ITL4=100 TRTOL=7

16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.001 1e-005 1e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2736 8525888 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 118
0 0
4.85009e-315 0 5.4086e-315 5.28841e-315 4.85009e-315 4.85009e-315
16 0
4 0.0003 5
1
18 115
0 8 0 0 1	0 10 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
