CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 452
7 5.000 V
7 5.000 V
3 GND
0 66 640 452
9437186 0
0
0
0
0
0
0
16
14 Logic Display~
6 555 44 0 1 3
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8953 0 0
0
0
9 Inverter~
13 10 271 0 2 21
0 2 3
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U1B
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 -33686019
65 0 0 0 6 2 1 0
1 U
4441 0 0
0
0
10 Ascii Key~
169 34 209 0 11 11
0 9 8 7 6 45 46 47 2 0
0 48
0
0 0 20528 0
0
0
0
0
0
0
0
0
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3618 0 0
0
0
2 +V
167 76 204 0 1 3
0 10
0
0 0 53488 0
3 10V
12 -2 33 6
0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
7 74LS164
127 485 271 0 12 25
0 10 6 3 10 48 49 50 51 25
21 17 13
0
0 0 12528 0
7 74LS164
-24 -51 25 -43
0
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 -33686019
65 0 0 512 1 1 0 0
1 U
5394 0 0
0
0
7 74LS164
127 367 271 0 12 25
0 10 7 3 10 52 53 54 55 26
22 18 14
0
0 0 12528 0
7 74LS164
-24 -51 25 -43
0
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 -33686019
65 0 0 512 1 1 0 0
1 U
7734 0 0
0
0
7 74LS164
127 246 271 0 12 25
0 10 8 3 10 56 57 58 59 27
23 19 15
0
0 0 12528 0
7 74LS164
-24 -51 25 -43
0
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 -33686019
65 0 0 512 1 1 0 0
1 U
9914 0 0
0
0
7 74LS164
127 126 271 0 12 25
0 10 9 3 10 60 61 62 63 28
24 20 16
0
0 0 12528 0
7 74LS164
-24 -51 25 -43
0
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 -33686019
65 0 0 512 1 1 0 0
1 U
3747 0 0
0
0
6 74LS85
106 494 111 0 14 29
0 36 35 34 33 13 14 15 16 64
11 65 66 5 67
0
0 0 12528 0
6 74LS85
-21 -51 21 -43
0
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 -33686019
65 0 0 512 1 1 0 0
1 U
3549 0 0
0
0
6 74LS85
106 384 111 0 14 29
0 40 39 38 37 17 18 19 20 68
4 69 70 11 71
0
0 0 12528 0
6 74LS85
-21 -51 21 -43
0
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 -33686019
65 0 0 512 1 1 0 0
1 U
7931 0 0
0
0
6 74LS85
106 274 111 0 14 29
0 29 30 31 32 21 22 23 24 72
12 73 74 4 75
0
0 0 12528 0
6 74LS85
-21 -51 21 -43
0
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 -33686019
65 0 0 512 1 1 0 0
1 U
9325 0 0
0
0
6 74LS85
106 164 111 0 14 29
0 44 43 42 41 25 26 27 28 76
77 78 79 12 80
0
0 0 12528 0
6 74LS85
-21 -51 21 -43
0
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 -33686019
65 0 0 512 1 1 0 0
1 U
8903 0 0
0
0
8 Hex Key~
166 444 31 0 11 11
0 33 34 35 36 0 0 0 0 0
2 50
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3834 0 0
0
0
8 Hex Key~
166 334 31 0 11 11
0 37 38 39 40 0 0 0 0 0
4 52
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3363 0 0
0
0
8 Hex Key~
166 224 31 0 11 11
0 32 31 30 29 0 0 0 0 0
7 55
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7668 0 0
0
0
8 Hex Key~
166 113 32 0 11 11
0 41 42 43 44 0 0 0 0 0
1 49
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4718 0 0
0
0
70
8 1 2 0 0 4224 0 3 2 0 0 2
13 233
13 253
2 3 3 0 0 8320 0 2 5 0 0 5
13 289
13 337
448 337
448 271
453 271
3 0 3 0 0 0 0 8 0 0 2 3
94 271
64 271
64 337
3 0 3 0 0 0 0 7 0 0 2 3
214 271
204 271
204 337
3 0 3 0 0 0 0 6 0 0 2 3
335 271
324 271
324 337
13 10 4 0 0 12416 0 11 10 0 0 6
306 138
315 138
315 61
420 61
420 93
416 93
1 13 5 0 0 4224 0 1 9 0 0 3
555 62
555 138
526 138
4 2 6 0 0 8320 0 3 5 0 0 5
37 233
37 331
441 331
441 253
453 253
3 2 7 0 0 8320 0 3 6 0 0 5
43 233
43 326
310 326
310 253
335 253
2 2 8 0 0 8320 0 3 7 0 0 5
49 233
49 320
190 320
190 253
214 253
2 1 9 0 0 4224 0 8 3 0 0 3
94 253
55 253
55 233
1 0 10 0 0 4096 0 8 0 0 13 2
94 244
76 244
4 0 10 0 0 8192 0 8 0 0 19 3
88 289
76 289
76 219
1 0 10 0 0 0 0 7 0 0 15 2
214 244
197 244
4 0 10 0 0 0 0 7 0 0 19 3
208 289
197 289
197 219
1 0 10 0 0 0 0 6 0 0 17 2
335 244
317 244
4 0 10 0 0 0 0 6 0 0 19 3
329 289
317 289
317 219
1 0 10 0 0 0 0 5 0 0 19 2
453 244
434 244
1 4 10 0 0 8320 0 4 5 0 0 5
76 213
76 219
434 219
434 289
447 289
13 10 11 0 0 12416 0 10 9 0 0 6
416 138
426 138
426 62
534 62
534 93
526 93
10 13 12 0 0 12416 0 11 12 0 0 6
306 93
310 93
310 62
204 62
204 138
196 138
12 16 13 0 0 8320 0 5 0 0 54 3
517 307
544 307
544 191
12 15 14 0 0 8320 0 6 0 0 54 3
399 307
427 307
427 191
12 14 15 0 0 8320 0 7 0 0 54 3
278 307
303 307
303 191
12 13 16 0 0 8320 0 8 0 0 54 3
158 307
183 307
183 191
11 12 17 0 0 8320 0 5 0 0 54 3
517 298
536 298
536 191
11 11 18 0 0 8320 0 6 0 0 54 3
399 298
419 298
419 191
11 10 19 0 0 8320 0 7 0 0 54 3
278 298
296 298
296 191
11 9 20 0 0 8320 0 8 0 0 54 3
158 298
176 298
176 191
10 8 21 0 0 8320 0 5 0 0 54 3
517 289
528 289
528 191
10 7 22 0 0 8320 0 6 0 0 54 3
399 289
410 289
410 191
10 6 23 0 0 8320 0 7 0 0 54 3
278 289
289 289
289 191
10 5 24 0 0 8320 0 8 0 0 54 3
158 289
168 289
168 191
9 4 25 0 0 8320 0 5 0 0 54 3
517 280
521 280
521 191
9 3 26 0 0 8320 0 6 0 0 54 3
399 280
402 280
402 191
9 2 27 0 0 8320 0 7 0 0 54 3
278 280
282 280
282 191
9 1 28 0 0 8320 0 8 0 0 54 3
158 280
161 280
161 191
5 16 13 0 0 0 0 9 0 0 54 3
462 120
431 120
431 191
6 15 14 0 0 0 0 9 0 0 54 3
462 129
439 129
439 191
7 14 15 0 0 0 0 9 0 0 54 3
462 138
448 138
448 191
8 13 16 0 0 0 0 9 0 0 54 3
462 147
456 147
456 191
5 12 17 0 0 0 0 10 0 0 54 3
352 120
320 120
320 191
6 11 18 0 0 0 0 10 0 0 54 3
352 129
329 129
329 191
7 10 19 0 0 0 0 10 0 0 54 3
352 138
337 138
337 191
8 9 20 0 0 0 0 10 0 0 54 3
352 147
344 147
344 191
5 8 21 0 0 0 0 11 0 0 54 3
242 120
211 120
211 191
6 7 22 0 0 0 0 11 0 0 54 3
242 129
219 129
219 191
7 6 23 0 0 0 0 11 0 0 54 3
242 138
226 138
226 191
8 5 24 0 0 0 0 11 0 0 54 3
242 147
233 147
233 191
5 4 25 0 0 0 0 12 0 0 54 3
132 120
100 120
100 191
6 3 26 0 0 0 0 12 0 0 54 3
132 129
108 129
108 191
7 2 27 0 0 0 0 12 0 0 54 3
132 138
116 138
116 191
8 1 28 0 0 0 0 12 0 0 54 3
132 147
123 147
123 191
1 0 1 0 0 4256 0 0 0 0 0 2
93 191
575 191
1 4 29 0 0 8320 0 11 15 0 0 3
242 84
215 84
215 55
3 2 30 0 0 4224 0 15 11 0 0 3
221 55
221 93
242 93
3 2 31 0 0 8320 0 11 15 0 0 3
242 102
227 102
227 55
1 4 32 0 0 4224 0 15 11 0 0 3
233 55
233 111
242 111
1 4 33 0 0 4224 0 13 9 0 0 3
453 55
453 111
462 111
2 3 34 0 0 4224 0 13 9 0 0 3
447 55
447 102
462 102
3 2 35 0 0 4224 0 13 9 0 0 3
441 55
441 93
462 93
4 1 36 0 0 4224 0 13 9 0 0 3
435 55
435 84
462 84
1 4 37 0 0 4224 0 14 10 0 0 3
343 55
343 111
352 111
2 3 38 0 0 4224 0 14 10 0 0 3
337 55
337 102
352 102
3 2 39 0 0 4224 0 14 10 0 0 3
331 55
331 93
352 93
4 1 40 0 0 4224 0 14 10 0 0 3
325 55
325 84
352 84
1 4 41 0 0 4224 0 16 12 0 0 3
122 56
122 111
132 111
2 3 42 0 0 4224 0 16 12 0 0 3
116 56
116 102
132 102
3 2 43 0 0 4224 0 16 12 0 0 3
110 56
110 93
132 93
4 1 44 0 0 4224 0 16 12 0 0 3
104 56
104 84
132 84
7
16 8 0 0 0 0 0 0 0 0 0 0 54
6 System
0 0 0 4
532 8 580 30
536 12 570 28
4 Open
16 8 0 0 0 0 0 0 0 0 0 0 54
6 System
0 0 0 25
3 5 98 46
7 9 88 41
25 Combination
Lock Circuit
16 8 0 0 0 0 0 0 0 0 0 0 54
6 System
0 0 0 12
129 5 177 46
133 9 167 41
12 First
Digit
16 8 0 0 0 0 0 0 0 0 0 0 54
6 System
0 0 0 13
239 6 301 47
243 10 291 42
13 Second
Digit
16 8 0 0 0 0 0 0 0 0 0 0 54
6 System
0 0 0 12
351 6 399 47
355 10 389 42
12 Third
Digit
16 8 0 0 0 0 0 0 0 0 0 0 54
6 System
0 0 0 13
459 5 514 46
463 9 504 41
13 Fourth
Digit
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 133
0 38 105 211
4 42 102 182
133 Click on the 
key symbol 
below to 
select it 
then press 
the correct 
digits on 
the keyboard 
to open the 
lock.
0
17 0 0
0
0
3 Vin
-1.5 -0.7 0.01
3 Vcc
10 14 1
100 0 1 100000
0 0.0005 2.5e-006 2.5e-006 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 100 100 0 0
77 66 617 126
0 0 0 0
617 66
77 66
617 66
617 126
0 0
1e-007 0 12 -12 1e-007 1e-007
16 0
0 3e-008 5
0
0 0 100 100 0 0
98 66 294 126
0 0 0 0
294 66
98 66
294 66
294 126
0 0
1e+007 1 12.16 12.184 1e+007 1e+007
12403 0
0 3e+006 5e+006
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
2000 1 2.38857 0 1999 1999
16 0
0 500 1000
0
0 0 100 100 0 0
98 66 296 126
0 0 0 0
296 66
98 66
296 66
296 126
0 0
1e+006 1 -3.55271e-015 0 999999 999999
12403 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
