CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
52 C:\Users\Jefferson\Desktop\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1446 465
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 142 403 0 1 11
0 10
0
0 0 21360 0
2 0V
-29 -4 -15 4
1 C
-4 -32 3 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7159 0 0
2
44111.9 0
0
13 Logic Switch~
5 146 192 0 1 11
0 7
0
0 0 21360 0
2 0V
-29 -4 -15 4
1 A
-4 -32 3 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5812 0 0
2
44111.9 0
0
13 Logic Switch~
5 143 301 0 1 11
0 8
0
0 0 21360 0
2 0V
-29 -4 -15 4
1 B
-4 -32 3 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
331 0 0
2
44111.9 0
0
8 4-In OR~
219 430 306 0 5 22
0 5 6 4 13 3
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 3 0
1 U
9604 0 0
2
44111.9 0
0
5 4073~
219 326 396 0 4 22
0 7 8 9 4
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
7518 0 0
2
44111.9 0
0
5 4073~
219 327 302 0 4 22
0 7 11 10 6
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
4832 0 0
2
44111.9 0
0
5 4073~
219 325 202 0 4 22
0 12 8 10 5
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
6798 0 0
2
44111.9 0
0
9 Inverter~
13 260 404 0 2 22
0 10 9
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3336 0 0
2
44111.9 1
0
9 Inverter~
13 264 193 0 2 22
0 7 12
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
8370 0 0
2
44111.9 1
0
9 Inverter~
13 261 302 0 2 22
0 8 11
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3910 0 0
2
44111.9 0
0
4 LED~
171 516 330 0 2 2
10 3 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
316 0 0
2
44111.9 0
0
7 Ground~
168 516 358 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
536 0 0
2
44111.9 0
0
17
5 1 3 0 0 4224 0 4 11 0 0 3
463 306
516 306
516 320
4 3 4 0 0 8320 0 5 4 0 0 4
347 396
354 396
354 311
413 311
4 1 5 0 0 8320 0 7 4 0 0 4
346 202
354 202
354 293
413 293
4 2 6 0 0 4224 0 6 4 0 0 2
348 302
413 302
1 0 7 0 0 8192 0 5 0 0 9 3
302 387
209 387
209 293
2 0 8 0 0 4096 0 5 0 0 16 3
302 396
201 396
201 302
2 3 9 0 0 8320 0 8 5 0 0 3
281 404
281 405
302 405
3 0 10 0 0 4096 0 6 0 0 14 3
303 311
192 311
192 404
1 0 7 0 0 4224 0 6 0 0 15 3
303 293
191 293
191 193
2 2 11 0 0 4224 0 10 6 0 0 2
282 302
303 302
0 3 10 0 0 4224 0 0 7 14 0 3
181 404
181 211
301 211
0 2 8 0 0 8320 0 0 7 16 0 3
168 302
168 202
301 202
2 1 12 0 0 4224 0 9 7 0 0 2
285 193
301 193
1 1 10 0 0 16 0 1 8 0 0 3
154 403
154 404
245 404
1 1 7 0 0 0 0 2 9 0 0 3
158 192
158 193
249 193
1 1 8 0 0 0 0 3 10 0 0 3
155 301
155 302
246 302
1 2 2 0 0 4224 0 12 11 0 0 4
516 352
516 339
516 339
516 340
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
