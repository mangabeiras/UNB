CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 9 100 3
0 70 640 452
7 5.000 V
7 5.000 V
3 GND
0 70 640 452
11534338 0
0
0
0
0
0
0
24
13 Logic Switch~
5 34 134 0 1 3
0 11
0
0 0 112 0
2 0V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 35 103 0 1 3
0 12
0
0 0 112 0
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 35 71 0 1 3
0 13
0
0 0 112 0
2 0V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 35 38 0 1 3
0 14
0
0 0 112 0
2 0V
-7 -16 7 -8
2 V4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Piezo Buzzer~
174 362 289 0 2 5
10 3 2
0
0 0 4208 0
4 .1uF
10 -16 38 -8
3 BZ1
13 -26 34 -18
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
2 BZ
5394 0 0
0
0
9 DC Motor~
219 369 223 0 2 5
0 5 2
0
0 0 112 0
4 100H
-15 -42 13 -34
2 M1
-8 -52 6 -44
0
0
27 %D %1 N%D %V
R%D N%D %2 10
0
0
0
5

0 0 0 0 0 0
76 0 0 0 0 0 0 0
1 M
7734 0 0
0
0
9 DC Motor~
219 367 63 0 2 5
0 10 2
0
0 0 112 0
4 100H
-15 -42 13 -34
2 M2
-8 -52 6 -44
0
0
27 %D %1 N%D %V
R%D N%D %2 10
0
0
0
5

0 0 0 0 0 0
76 0 0 0 0 0 0 0
1 M
9914 0 0
0
0
13 Relay Coil:A~
209 371 168 0 2 5
0 6 2
0
0 0 5232 90
8 120VCOIL
-28 -44 28 -36
4 RLY1
-14 -54 14 -46
2 K1
-10 -24 4 -16
0
24 *p=1 r=1
%D %1 %2 %I %S
0
39 alias:XCOIL {PULLIN=96 RESISTANCE=2000}
0
5

0 1 2 1 2 0
88 0 0 0 0 0 -2 0
3 RLY
3747 0 0
0
0
11 Contacts:D~
214 247 222 0 3 7
0 5 15 4
0
0 0 17520 0
6 NORMAL
-21 -44 21 -36
4 RLY2
-14 -54 14 -46
2 K1
-6 -20 8 -12
0
18 %D %1 %3 N%D %I %S
0
15 alias:XCONTACTS
0
7

0 1 2 3 1 2 3 0
88 0 0 0 0 0 -2 0
3 RLY
3549 0 0
0
0
9 Solenoid~
210 88 134 0 2 5
0 11 2
0
0 0 5232 0
6 5VCOIL
-21 -44 21 -36
4 RLY3
-14 -54 14 -46
2 S4
-7 -16 7 -8
0
24 *p=1 r=1
%D %1 %2 %I %S
0
11 alias:XCOIL
0
5

0 1 2 1 2 0
88 0 0 0 0 0 -3 0
3 RLY
7931 0 0
0
0
9 Solenoid~
210 86 103 0 2 5
0 12 2
0
0 0 5232 0
6 5VCOIL
-21 -44 21 -36
4 RLY4
-14 -54 14 -46
2 S3
-7 -16 7 -8
0
24 *p=1 r=1
%D %1 %2 %I %S
0
11 alias:XCOIL
0
5

0 1 2 1 2 0
88 0 0 0 0 0 -4 0
3 RLY
9325 0 0
0
0
9 Solenoid~
210 87 71 0 2 5
0 13 2
0
0 0 5232 0
6 5VCOIL
-21 -44 21 -36
4 RLY5
-14 -54 14 -46
2 S2
-7 -16 7 -8
0
24 *p=1 r=1
%D %1 %2 %I %S
0
11 alias:XCOIL
0
5

0 1 2 1 2 0
88 0 0 0 0 0 -5 0
3 RLY
8903 0 0
0
0
11 Contacts:D~
214 311 131 0 3 7
0 7 16 4
0
0 0 17520 0
6 NORMAL
-21 -44 21 -36
4 RLY6
-14 -54 14 -46
2 S4
-6 -20 8 -12
0
18 %D %1 %3 N%D %I %S
0
15 alias:XCONTACTS
0
7

0 1 2 3 1 2 3 0
88 0 0 0 0 0 -3 0
3 RLY
3834 0 0
0
0
11 Contacts:D~
214 312 62 0 3 7
0 10 17 8
0
0 0 17520 0
6 NORMAL
-21 -44 21 -36
4 RLY7
-14 -54 14 -46
2 S4
-6 -19 8 -11
0
18 %D %1 %3 N%D %I %S
0
15 alias:XCONTACTS
0
7

0 1 2 3 1 2 3 0
88 0 0 0 0 0 -3 0
3 RLY
3363 0 0
0
0
11 Contacts:D~
214 234 93 0 3 7
0 8 18 4
0
0 0 17520 0
6 NORMAL
-21 -44 21 -36
4 RLY8
-14 -54 14 -46
2 S3
-6 -19 8 -11
0
18 %D %1 %3 N%D %I %S
0
15 alias:XCONTACTS
0
7

0 1 2 3 1 2 3 0
88 0 0 0 0 0 -4 0
3 RLY
7668 0 0
0
0
11 Contacts:D~
214 213 62 0 3 7
0 8 19 4
0
0 0 17520 0
6 NORMAL
-21 -44 21 -36
4 RLY9
-14 -54 14 -46
2 S1
-7 -20 7 -12
0
18 %D %1 %3 N%D %I %S
0
15 alias:XCONTACTS
0
7

0 1 2 3 1 2 3 0
88 0 0 0 0 0 -6 0
3 RLY
4718 0 0
0
0
9 Solenoid~
210 88 38 0 2 5
0 14 2
0
0 0 5232 0
6 5VCOIL
-21 -44 21 -36
5 RLY10
-18 -54 17 -46
2 S1
-7 -16 7 -8
0
24 *p=1 r=1
%D %1 %2 %I %S
0
11 alias:XCOIL
0
5

0 1 2 1 2 0
88 0 0 0 0 0 -6 0
3 RLY
3874 0 0
0
0
11 Contacts:E~
214 259 62 0 3 7
0 8 8 20
0
0 0 17520 0
6 NORMAL
-21 -44 21 -36
5 RLY11
-18 -54 17 -46
2 S2
-6 -21 8 -13
0
18 %D %1 N%D %2 %I %S
0
15 alias:XCONTACTS
0
7

0 1 2 3 1 2 3 0
88 0 0 0 0 0 -5 0
3 RLY
6671 0 0
0
0
14 NO PushButton~
191 250 281 0 2 5
0 3 4
0
0 0 20592 0
0
2 S1
-7 -30 7 -22
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3789 0 0
0
0
14 NO PushButton~
191 249 179 0 2 5
0 6 4
0
0 0 20592 0
0
2 S2
-7 -30 7 -22
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
4871 0 0
0
0
5 Lamp~
206 369 118 0 2 5
11 7 2
0
0 0 96 0
3 100
-10 -24 11 -16
2 L1
-7 -34 7 -26
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3750 0 0
0
0
7 Ground~
168 406 325 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8778 0 0
0
0
2 +V
167 181 37 0 1 3
0 4
0
0 0 53488 0
3 10V
12 -2 33 6
2 V5
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
538 0 0
0
0
7 Ground~
168 128 156 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
2

0 1 0
0 0 0 0 1 0 0 0
0
6843 0 0
0
0
29
2 0 2 0 0 4096 0 5 0 0 20 2
393 289
406 289
1 1 3 0 0 4224 0 19 5 0 0 2
267 289
331 289
2 0 4 0 0 4096 0 19 0 0 21 2
233 289
181 289
2 0 2 0 0 0 0 6 0 0 20 2
393 222
406 222
1 1 5 0 0 4224 0 9 6 0 0 2
265 222
345 222
3 0 4 0 0 0 0 9 0 0 21 2
229 222
181 222
2 0 2 0 0 8192 0 8 0 0 20 3
380 181
380 186
406 186
1 1 6 0 0 4224 0 20 8 0 0 3
266 187
356 187
356 181
2 0 4 0 0 0 0 20 0 0 21 2
232 187
181 187
2 0 2 0 0 0 0 21 0 0 20 2
381 131
406 131
1 1 7 0 0 4224 0 13 21 0 0 2
329 131
357 131
3 0 4 0 0 4096 0 13 0 0 21 2
293 131
181 131
1 0 8 0 0 4224 0 15 0 0 17 3
252 93
286 93
286 62
3 0 4 0 0 0 0 15 0 0 21 2
216 93
181 93
3 0 4 0 0 0 0 16 0 0 21 2
195 62
181 62
2 1 8 0 0 4224 9 18 16 0 0 2
241 62
231 62
3 1 8 0 0 0 0 14 18 0 0 2
294 62
277 62
1 1 10 0 0 4224 0 7 14 0 0 2
343 62
330 62
2 0 2 0 0 0 0 7 0 0 20 2
391 62
406 62
1 0 2 0 0 4224 0 22 0 0 0 2
406 319
406 27
1 0 4 0 0 4224 0 23 0 0 0 2
181 46
181 333
2 0 2 0 0 0 0 10 0 0 25 2
108 134
128 134
2 0 2 0 0 0 0 11 0 0 25 2
106 103
128 103
2 0 2 0 0 0 0 12 0 0 25 2
107 71
128 71
2 1 2 0 0 0 0 17 24 0 0 3
108 38
128 38
128 150
1 1 11 0 0 4224 0 1 10 0 0 2
46 134
68 134
1 1 12 0 0 4224 0 2 11 0 0 2
47 103
66 103
1 1 13 0 0 4224 0 3 12 0 0 2
47 71
67 71
1 1 14 0 0 4224 0 4 17 0 0 2
47 38
68 38
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 2e-006 1e-008 1e-008 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
3524 1210432 100 100 0 0
0 0 0 0
0 66 140 136
0 0
0 0
0 0
0 0
0 0
5.43943e-315 5.2221e-315 5.5705e-315 0 5.43813e-315 5.5705e-315
16 0
4 1 100
1
339 131
0 7 0 0 1	0 11 0 0
1120 8550464 100 100 0 0
77 66 617 126
14 477 654 670
617 66
77 66
617 66
617 126
0 0
4.78936e-315 0 5.27018e-315 5.10937e-315 4.80864e-315 4.80864e-315
16 0
4 5e-007 100
1
330 62
0 10 0 0 1	0 18 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
