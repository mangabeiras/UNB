CircuitMaker Text
5.6
Probes: 6
U1_6
Fourier Analysis
0 199 70 65280
out
Operating Point
0 198 65 65280
out
DC Sweep
0 198 67 65280
out
AC Analysis
0 198 67 65280
out
Transient Analysis
0 198 67 65280
Vin_1
Transient Analysis
1 76 87 65535
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 10
245 80 857 634
7 5.000 V
7 5.000 V
3 GND
10000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
2 4 0.500000 0.500000
413 176 1025 453
12058632 0
0
0
0
0
0
0
9
7 Ground~
168 198 158 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
5130 0 0
2
36626.4 1
0
2 +V
167 153 135 0 1 64
0 5
0
0 0 54128 180
4 -12V
-14 0 14 8
3 Vee
-9 10 12 18
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
391 0 0
2
36626.4 2
0
2 +V
167 153 59 0 1 64
0 4
0
0 0 54128 0
4 +12v
-13 -13 15 -5
3 Vcc
-9 -23 12 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
36626.4 3
0
7 Ground~
168 101 131 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3421 0 0
2
36626.4 4
0
11 Signal Gen~
195 41 93 0 19 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 -1110651699 1176256512 0 1036831949
20
-0.1 10000 0 0.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -100m/100mV
-38 23 39 31
3 Vin
-11 -31 10 -23
0
0
44 %D %1 %2 DC 0 SIN(0 100m 10k 0 0) AC -100m 0
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
36626.4 5
0
8 Op-Amp5~
219 153 94 0 5 64
0 2 6 4 5 3
8 Op-Amp5~
0 0 848 0
5 UA741
7 -13 42 -5
2 U1
15 -23 29 -15
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 -33686019
88 0 0 0 1 0 0 0
1 U
5572 0 0
2
36626.4 6
0
9 Resistor~
219 101 88 0 2 64
0 7 6
9 Resistor~
0 0 4976 0
3 10k
-10 -12 11 -4
2 RI
-6 -23 8 -15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8901 0 0
2
36626.4 7
0
9 Resistor~
219 164 25 0 2 64
0 6 3
9 Resistor~
0 0 4976 0
6 100.0k
-20 -12 22 -4
2 RF
-6 -22 8 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7361 0 0
2
36626.4 8
0
9 Resistor~
219 198 122 0 3 64
0 2 3 -1
9 Resistor~
0 0 4976 90
3 25k
5 1 26 9
2 RL
7 -9 21 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4747 0 0
2
36626.4 9
0
10
1 0 2 0 0 4096 0 4 0 0 2 2
101 125
101 100
1 2 2 0 0 4224 0 6 5 0 0 4
135 100
83 100
83 98
72 98
1 1 2 0 0 0 0 9 1 0 0 2
198 140
198 152
3 1 4 0 0 4224 0 6 3 0 0 2
153 81
153 68
4 1 5 0 0 4224 0 6 2 0 0 2
153 107
153 120
1 0 6 0 0 8320 0 8 0 0 7 3
146 25
127 25
127 88
2 2 6 0 0 0 0 7 6 0 0 2
119 88
135 88
2 0 3 0 0 8320 0 8 0 0 9 3
182 25
198 25
198 94
5 2 3 0 0 0 0 6 9 0 0 3
171 94
198 94
198 104
1 1 7 0 0 4224 0 5 7 0 0 2
72 88
83 88
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 3
198 46 225 62
198 46 225 62
3 out
0
29 0 1
0
0
3 Vin
-0.7 -1.5 -0.02
0
0 0 0
100 0 1 1e+06
0 0.0005 2.5e-06 2.5e-06
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3236 1210432 100 100 0 0
77 66 617 126
0 66 140 136
617 66
77 66
617 66
617 126
0 0
0 0 0 0 0 0
16 0
4 1 5
1
153 76
0 3 0 0 1	0 4 0 0
756 8550464 100 100 0 0
77 66 287 126
0 259 320 452
286 66
77 66
287 66
287 126
0 0
0 0 0 0 0 0
16 0
4 0.0001 5
2
78 88
0 7 0 0 1	0 10 0 0
198 60
0 6 0 0 2	0 8 0 0
3552 2259008 100 100 0 0
77 66 287 126
320 66 640 259
287 66
77 66
287 66
287 126
0 0
0 0 0 0 0 0
0 0
4 0.3 5
1
198 62
0 6 0 0 2	0 8 0 0
3600 4421696 100 100 0 0
98 66 296 126
320 259 640 452
296 66
98 66
296 66
296 66
0 0
0 0 0 0 0 0
12403 0
4 300000 500000
1
198 67
0 6 0 0 2	0 8 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
