CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 507 352
7 5.000 V
7 5.000 V
3 GND
1666.67 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 507 352
9961474 0
0
0
0
0
0
0
12
5 SAVE-
218 413 59 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
26 *Combine
*TRAN -17m 17.3m
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 72 66 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
26 *Combine
*TRAN -17m 17.3m
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
11 Signal Gen~
195 41 91 0 19 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 981668463
20
1 1000 0 0.001 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 576 0
5 -1/1V
-15 -48 20 -40
2 V1
-8 -30 6 -22
0
0
37 %D %1 %2 DC 0 SIN(0 1m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
7 Ground~
168 221 173 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
8 Battery~
219 149 129 0 2 64
0 2 7
8 Battery~
0 0 832 180
2 5V
-29 -3 -15 5
2 V2
-29 -13 -15 -5
0
0
14 %D %1 %2 DC %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 1 0 0
1 V
5394 0 0
0
0
10 NPN Trans~
219 222 38 0 3 64
0 4 2 3
10 NPN Trans~
0 0 832 602
6 2N3904
-19 -18 23 -10
2 Q1
-4 -30 10 -22
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 0 0 0 1 0 0 0
1 Q
7734 0 0
0
0
8 Battery~
219 309 124 0 2 64
0 8 2
8 Battery~
0 0 832 0
3 12V
11 -3 32 5
2 V3
15 -14 29 -6
0
0
14 %D %1 %2 DC %V
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 1 0 0
1 V
9914 0 0
0
0
10 Polar Cap~
219 113 30 0 2 64
0 6 3
10 Polar Cap~
0 0 832 0
3 1uF
-12 -18 9 -10
2 C1
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
10 Polar Cap~
219 375 30 0 2 64
0 4 5
10 Polar Cap~
0 0 832 0
3 1uF
-12 -18 9 -10
2 C2
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
9 Resistor~
219 309 75 0 2 64
0 8 4
9 Resistor~
0 0 4960 90
4 4.7K
5 -1 33 7
2 R1
7 -12 21 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 147 73 0 2 64
0 7 3
9 Resistor~
0 0 4960 90
4 4.7K
6 -1 34 7
2 R2
7 -12 21 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 413 91 0 3 64
0 2 5 -1
9 Resistor~
0 0 4960 90
3 10K
6 -1 27 7
2 R3
12 -11 26 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
13
2 0 2 0 0 4096 0 6 0 0 10 2
221 43
221 156
3 2 3 0 0 4224 0 6 11 0 0 3
203 30
147 30
147 55
1 2 4 0 0 4224 0 6 10 0 0 3
239 30
309 30
309 57
1 0 2 0 0 0 0 12 0 0 11 3
413 109
413 156
309 156
2 2 5 0 0 8320 0 9 12 0 0 3
381 30
413 30
413 73
0 1 4 0 0 0 0 0 9 3 0 2
309 30
364 30
2 0 2 0 0 0 0 3 0 0 11 3
72 96
72 156
147 156
1 1 6 0 0 8320 0 8 3 0 0 3
102 30
72 30
72 86
2 0 3 0 0 0 0 8 0 0 2 2
119 30
147 30
1 0 2 0 0 0 0 4 0 0 11 2
221 167
221 156
1 2 2 0 0 8320 0 5 7 0 0 4
147 138
147 156
309 156
309 135
2 1 7 0 0 4224 0 5 11 0 0 2
147 114
147 91
1 1 8 0 0 4224 0 7 10 0 0 2
309 111
309 93
0
0
16 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.003 1e-005 1e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1120 8550464 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
0 0 0 0 0 0
16 0
4 0.001 5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
