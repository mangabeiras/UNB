CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 20 9
0 66 640 452
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 452
11534336 0
1
19 2 Channel Audio Amp
12 John Adamson
7 9-18-93
7 12-7-94
18 Not for Simulation
207
4 LED~
171 685 32 0 64 64
10 2 9 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
0
0 0 17008 90
4 LED0
-12 -21 16 -13
4 LED3
-12 -24 16 -16
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8953 0 0
0
0
2 +V
167 829 22 0 64 64
0 10 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
0
0 0 53600 0
4 -30V
-13 -14 15 -6
3 V12
-10 -24 11 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
7 Output~
178 856 53 0 64 64
0 3 0 0 0 0 0 0 0 0
67 104 50 32 68 105 114 32 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
0
0 0 53344 0
0
0
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3618 0 0
0
0
12 SPDT Switch~
164 791 37 0 3 11
0 10 8 116
0
0 0 20832 -757982208
2 S1
-7 -17 7 -9
2 S1
-7 -27 7 -19
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 -1 0
1 S
6153 0 0
0
0
12 SPDT Switch~
164 791 53 0 3 11
0 3 11 117
0
0 0 20576 -757982208
2 S1
-7 -15 7 -7
2 S2
-7 -25 7 -17
0
0
0
0
0
0
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 -1 0
1 S
5394 0 0
0
0
7 Ground~
168 649 103 0 64 64
0 2 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
5 Coax~
219 703 82 0 64 64
0 7 2 11 118 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
5 Coax~
0 0 16640 0
12 Coax Cable 3
-42 -20 42 -12
5 CABL1
-18 -30 17 -22
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 252 512 1 0 0 0
4 CABL
9914 0 0
0
0
2 +V
167 2210 274 0 1 64
0 13
0
0 0 53600 23685390
4 +15V
8 -5 36 3
2 V1
15 -15 29 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
2 +V
167 2166 79 0 1 64
0 16
0
0 0 53600 0
4 +15V
-13 -13 15 -5
2 V2
-6 -23 8 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
2 +V
167 2120 64 0 1 64
0 17
0
0 0 53600 0
4 -15V
-15 -13 13 -5
2 V3
-8 -23 6 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
7 Ground~
168 1998 288 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
7 Ground~
168 2262 72 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
12 SPST Switch~
165 2314 86 0 2 11
0 2 20
0
0 0 21088 90
0
3 TC1
-32 -5 -11 3
0
0
0
0
0
0
5

0 1 2 1 2 -33686019
0 0 0 0 1 0 0 0
1 S
3834 0 0
0
0
6 Diode~
219 2280 229 0 2 64
0 20 23
6 Diode~
0 0 832 46260
6 1N4002
-21 -18 21 -10
3 D13
-11 -28 10 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 -1 280 0 1 0 0 0
1 D
3363 0 0
0
0
8 Op-Amp5~
219 2166 132 0 5 64
0 14 18 16 119 22
8 Op-Amp5~
0 0 832 0
5 LM358
7 -15 42 -7
3 U1A
14 -25 35 -17
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
64

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 255198399 141460666 439812096 77
459752504 145780 11010060 206045352 -2065956862 343 2097152 3933184 2228518 3670334
-2068184920 1144546382 145780 134216 224330071 -2065038466 398426855 0 5052983 41681930
9043980 34072 41817815 6079 439812096 67764301 385294670 439812096 923960600 439812096
77 41681930 25756284 77 6747516 76 -1070202874 6747516 385297432 -1074326058
335 6747432 343 -1074325948 9096152
88 -1 258 512 2 1 2 0
1 U
7668 0 0
0
0
8 Op-Amp5~
219 2166 229 0 5 64
0 15 14 120 121 24
8 Op-Amp5~
0 0 832 0
5 LM358
8 -13 43 -5
3 U1B
15 -23 36 -15
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
64

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 255198399 141460666 439812096 77
459752504 145780 11010060 206045352 -2065956862 343 2097152 3933184 2228518 3670334
-2068184920 1144546382 145780 134216 224330071 -2065038466 398426855 0 5052983 41681930
9043980 34072 41817815 6079 439812096 67764301 385294670 439812096 923960600 439812096
77 41681930 25756284 77 6747516 76 -1070202874 6747516 385297432 -1074326058
335 6747432 343 -1074325948 9096152
88 -1 258 512 2 2 2 0
1 U
4718 0 0
0
0
6 Diode~
219 2279 132 0 2 64
0 20 21
6 Diode~
0 0 832 46260
6 1N4002
-21 -18 21 -10
3 D12
-11 -28 10 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 -1 280 0 1 0 0 0
1 D
3874 0 0
0
0
7 Ground~
168 2028 681 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
7 Ground~
168 1966 681 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
3789 0 0
0
0
2 +V
167 2118 621 0 1 64
0 27
0
0 0 53600 23685390
4 -Vcc
6 -5 34 3
0
0
0
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
1 V
4871 0 0
0
0
5 Fuse~
219 2071 620 0 2 64
0 26 27
5 Fuse~
0 0 4928 0
3 10A
-10 -16 11 -8
2 F2
-7 -26 7 -18
0
0
11 %D %1 %2 %S
0
0
4 FUSE
5

0 1 2 1 2 -33686019
88 0 246 0 1 0 0 0
1 F
3750 0 0
0
0
2 +V
167 2041 43 0 1 64
0 28
0
0 0 53600 23685390
4 +Vcc
6 -5 34 3
0
0
0
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
1 V
8778 0 0
0
0
9 Terminal~
194 1973 352 0 1 64
0 4
0
0 0 20736 23685390
6 Output
6 -5 48 3
2 T1
20 -15 34 -7
0
0
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
1 T
538 0 0
0
0
7 Ground~
168 1905 470 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
6843 0 0
0
0
4 LED~
171 1871 397 0 2 64
10 31 30
0
0 0 624 90
4 LED0
-12 -21 16 -13
4 LED2
-10 13 18 21
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 -33686019
68 0 0 0 1 0 0 0
1 D
3136 0 0
0
0
7 Ground~
168 1799 513 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
2 +V
167 1780 338 0 1 64
0 32
0
0 0 53600 0
4 +12V
-14 -14 14 -6
2 V4
-7 -24 7 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
5670 0 0
0
0
11 SPDT Relay~
176 1835 362 0 10 64
0 29 122 4 32 31 0 0 0 0
1
0
0 0 21088 0
7 12VSPDT
-27 -35 22 -27
3 RY1
15 0 36 8
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 1 2 3 4 5 1 2 3 4
5 -33686019
88 0 0 512 1 0 0 0
3 RLY
6828 0 0
0
0
12 P-EMOS 3T:A~
219 1939 87 0 3 64
0 25 35 33
12 P-EMOS 3T:A~
0 0 832 46772
8 IRFP9240
13 12 69 20
3 Q19
28 1 49 9
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
109 0 552 0 1 0 0 0
1 Q
6735 0 0
0
0
12 P-EMOS 3T:A~
219 1820 87 0 3 64
0 25 36 33
12 P-EMOS 3T:A~
0 0 832 46772
8 IRFP9240
13 12 69 20
3 Q18
28 1 49 9
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
109 0 552 0 1 0 0 0
1 Q
8365 0 0
0
0
12 P-EMOS 3T:A~
219 1700 87 0 3 64
0 25 37 33
12 P-EMOS 3T:A~
0 0 832 46772
8 IRFP9240
13 12 69 20
3 Q17
28 1 49 9
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
109 0 552 0 1 0 0 0
1 Q
4132 0 0
0
0
12 N-EMOS 3T:A~
219 1939 596 0 3 64
0 25 39 26
12 N-EMOS 3T:A~
0 0 832 0
7 IRFP240
17 0 66 8
3 Q23
31 -10 52 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
77 0 546 0 1 0 0 0
1 Q
4551 0 0
0
0
12 N-EMOS 3T:A~
219 1820 596 0 3 64
0 25 40 26
12 N-EMOS 3T:A~
0 0 832 0
7 IRFP240
17 0 66 8
3 Q22
31 -10 52 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
77 0 546 0 1 0 0 0
1 Q
3635 0 0
0
0
12 N-EMOS 3T:A~
219 1700 597 0 3 64
0 25 41 26
12 N-EMOS 3T:A~
0 0 832 0
7 IRFP240
17 0 66 8
3 Q21
31 -10 52 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
77 0 546 0 1 0 0 0
1 Q
3973 0 0
0
0
12 Zener Diode~
219 1469 131 0 2 64
0 34 33
12 Zener Diode~
0 0 832 90
7 1N4742A
13 2 62 10
2 D6
31 -9 45 -1
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
100 0 281 0 1 0 0 0
1 D
3851 0 0
0
0
7 Ground~
168 1590 493 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
8383 0 0
0
0
2 +V
167 1494 502 0 1 64
0 46
0
0 0 53600 46260
4 +15V
-13 0 15 8
2 V5
-6 -10 8 -2
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
9334 0 0
0
0
2 +V
167 1494 414 0 1 64
0 47
0
0 0 53600 0
4 -15V
-13 -14 15 -6
2 V6
-6 -24 8 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
7471 0 0
0
0
7 Ground~
168 1353 368 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
3334 0 0
0
0
7 Ground~
168 1452 523 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
3559 0 0
0
0
12 PNP Trans:C~
219 1397 578 0 3 64
0 26 51 38
12 PNP Trans:C~
0 0 832 46772
6 MPSA56
18 0 60 8
3 Q15
29 -10 50 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
113 0 262 0 1 0 0 0
1 Q
984 0 0
0
0
4 LED~
171 1380 680 0 2 64
10 52 56
0
0 0 624 0
4 LED0
17 -5 45 3
4 LED1
18 -3 46 5
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 -33686019
68 0 0 0 1 0 0 0
1 D
7557 0 0
0
0
2 +V
167 1321 648 0 1 64
0 52
0
0 0 53600 0
4 +15V
-14 -14 14 -6
2 V7
-7 -24 7 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3146 0 0
0
0
7 Ground~
168 1321 812 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
5687 0 0
0
0
8 Caution~
219 850 815 0 1 64
0 0
8 Caution~
0 0 49248 0
0
0
0
0
0
0
0
0
3

0 0 0 -33686019
0 0 721 0 1 0 0 0
3 SYM
7939 0 0
0
0
11 Regulator3~
219 1100 629 0 3 64
0 59 58 57
11 Regulator3~
0 0 4864 0
6 LM337M
-21 -28 21 -20
3 IC9
-11 -38 10 -30
0
0
0
0
0
6 TO-220
7

0 3 1 2 3 1 2 -33686019
88 0 238 0 1 0 0 0
2 IC
3308 0 0
0
0
12 PNP Trans:C~
219 1329 557 0 3 64
0 51 61 62
12 PNP Trans:C~
0 0 832 46772
6 MPSA56
18 0 60 8
3 Q13
29 -10 50 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
113 0 262 0 1 0 0 0
1 Q
3408 0 0
0
0
12 PNP Trans:C~
219 1329 512 0 3 64
0 62 67 63
12 PNP Trans:C~
0 0 832 46772
6 MPSA56
18 0 60 8
3 Q12
29 -10 50 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
113 0 262 0 1 0 0 0
1 Q
9773 0 0
0
0
7 Ground~
168 1132 406 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
691 0 0
0
0
6 Diode~
219 1040 491 0 2 64
0 67 68
6 Diode~
0 0 832 90
6 1N4002
12 0 54 8
2 D2
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 -1 280 0 1 0 0 0
1 D
7834 0 0
0
0
12 Zener Diode~
219 1040 461 0 2 64
0 65 68
12 Zener Diode~
0 0 832 23685390
6 1N4728
14 -2 56 6
2 D4
28 -12 42 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
100 0 281 0 1 0 0 0
1 D
3588 0 0
0
0
12 NPN Trans:C~
219 1106 436 0 3 64
0 66 65 2
12 NPN Trans:C~
0 0 832 692
6 MPSA06
18 0 60 8
2 Q8
31 -10 45 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 -1 261 0 1 0 0 0
1 Q
4528 0 0
0
0
7 Ground~
168 1246 269 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
3303 0 0
0
0
7 Ground~
168 1402 188 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
9654 0 0
0
0
12 NPN Trans:C~
219 1329 246 0 3 64
0 70 73 64
12 NPN Trans:C~
0 0 832 0
6 MPSA06
18 0 60 8
3 Q11
28 -10 49 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 -1 261 0 1 0 0 0
1 Q
9791 0 0
0
0
12 NPN Trans:C~
219 1397 103 0 3 64
0 33 71 69
12 NPN Trans:C~
0 0 832 0
6 MPSA06
18 0 60 8
3 Q14
28 -10 49 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 -1 261 0 1 0 0 0
1 Q
4589 0 0
0
0
12 NPN Trans:C~
219 1329 137 0 3 64
0 71 80 70
12 NPN Trans:C~
0 0 832 0
6 MPSA06
18 0 60 8
3 Q10
28 -10 49 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 -1 261 0 1 0 0 0
1 Q
964 0 0
0
0
12 NPN Trans:C~
219 1263 295 0 3 64
0 66 72 2
12 NPN Trans:C~
0 0 832 692
6 MPSA06
18 0 60 8
2 Q9
31 -10 45 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 -1 261 0 1 0 0 0
1 Q
9151 0 0
0
0
2 +V
167 1175 361 0 1 64
0 74
0
0 0 53600 90
4 +15V
-33 -6 -5 2
2 V8
-26 -16 -12 -8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
4745 0 0
0
0
12 Zener Diode~
219 1176 295 0 2 64
0 77 76
12 Zener Diode~
0 0 832 0
6 1N4740
-21 -22 21 -14
2 D9
-7 -32 7 -24
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
100 0 281 0 1 0 0 0
1 D
8433 0 0
0
0
7 Ground~
168 1111 365 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
4221 0 0
0
0
12 NPN Trans:C~
219 1106 318 0 3 64
0 2 78 77
12 NPN Trans:C~
0 0 832 692
6 MPSA06
18 0 60 8
2 Q1
31 -10 45 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 -1 261 0 1 0 0 0
1 Q
8348 0 0
0
0
6 Diode~
219 1034 267 0 2 64
0 79 73
6 Diode~
0 0 832 90
6 1N4002
12 0 54 8
2 D1
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 -1 280 0 1 0 0 0
1 D
5299 0 0
0
0
12 Zener Diode~
219 1034 294 0 2 64
0 79 78
12 Zener Diode~
0 0 832 23685390
6 1N4728
14 -2 56 6
2 D3
28 -12 42 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
100 0 281 0 1 0 0 0
1 D
7393 0 0
0
0
2 +V
167 1111 227 0 1 64
0 75
0
0 0 53600 0
4 -15V
-14 -13 14 -5
2 V9
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
6917 0 0
0
0
7 Ground~
168 1212 113 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
8767 0 0
0
0
10 Capacitor~
219 1212 71 0 2 64
0 2 33
10 Capacitor~
0 0 832 90
5 100uF
11 0 46 8
3 C13
18 -10 39 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
3606 0 0
0
0
10 Capacitor~
219 1148 71 0 2 64
0 2 33
10 Capacitor~
0 0 832 90
4 .1uF
12 0 40 8
3 C12
15 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
6970 0 0
0
0
7 Ground~
168 877 296 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
343 0 0
0
0
12 NPN Trans:C~
219 931 541 0 3 64
0 67 87 86
12 NPN Trans:C~
0 0 832 0
6 MPSA06
18 0 60 8
2 Q6
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 -1 261 0 1 0 0 0
1 Q
7197 0 0
0
0
7 Ground~
168 625 665 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
3623 0 0
0
0
10 Capacitor~
219 625 638 0 2 64
0 2 59
10 Capacitor~
0 0 832 90
5 100uF
11 0 46 8
2 C3
22 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
7656 0 0
0
0
2 +V
167 598 622 0 1 64
0 59
0
0 0 53600 90
4 -30V
-35 -5 -7 3
3 V10
-32 -15 -11 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
5365 0 0
0
0
12 PNP Trans:C~
219 931 211 0 3 64
0 73 89 88
12 PNP Trans:C~
0 0 832 46772
6 MPSA56
18 0 60 8
2 Q5
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
113 0 262 0 1 0 0 0
1 Q
4557 0 0
0
0
7 Ground~
168 615 193 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
3489 0 0
0
0
2 +V
167 598 139 0 1 64
0 83
0
0 0 53600 90
4 +30V
-35 -5 -7 3
3 V11
-32 -15 -11 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
345 0 0
0
0
11 Regulator3~
219 716 409 0 3 64
0 83 95 94
11 Regulator3~
0 0 832 23685390
5 LM334
-15 -8 20 0
3 IC2
-8 -17 13 -9
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
88 0 238 0 1 1 0 0
1 U
3374 0 0
0
0
12 NPN Trans:C~
219 795 248 0 3 64
0 91 48 99
12 NPN Trans:C~
0 0 832 512
6 MPSA06
-64 0 -22 8
2 Q2
-50 -10 -36 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 -1 261 0 1 0 0 0
1 Q
5866 0 0
0
0
7 Ground~
168 641 55 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
631 0 0
0
0
10 Capacitor~
219 498 180 0 2 64
0 2 102
10 Capacitor~
0 0 832 0
5 .01uF
-18 -18 17 -10
3 C22
-11 -28 10 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
745 0 0
0
0
7 Ground~
168 477 279 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
7222 0 0
0
0
2 +V
167 519 147 0 1 64
0 102
0
0 0 53600 0
4 +15V
-13 -15 15 -7
3 V13
-10 -25 11 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
4508 0 0
0
0
8 Op-Amp5~
219 519 208 0 5 64
0 2 101 102 103 7
8 Op-Amp5~
0 0 832 0
5 LF357
12 18 47 26
3 IC6
19 6 40 14
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 -33686019
88 -1 258 0 1 0 0 0
1 U
3738 0 0
0
0
2 +V
167 519 287 0 1 64
0 103
0
0 0 53600 46260
4 -15V
-13 2 15 10
3 V14
-10 -8 11 0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
91 0 0
0
0
7 Ground~
168 543 446 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
4965 0 0
0
0
10 Capacitor~
219 487 374 0 2 64
0 104 106
10 Capacitor~
0 0 832 0
4 10uF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
7791 0 0
0
0
10 Capacitor~
219 571 400 0 2 64
0 2 105
10 Capacitor~
0 0 832 90
5 150pF
11 0 46 8
2 C2
22 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
3467 0 0
0
0
7 Ground~
168 427 386 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
3907 0 0
0
0
5 Coax~
219 434 315 0 4 64
0 107 123 104 2
5 Coax~
0 0 16640 270
12 Coax Cable 1
-95 7 -11 15
5 CABL2
-71 -3 -36 5
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -33686019
0 0 252 512 1 0 0 0
4 CABL
7505 0 0
0
0
9 Terminal~
194 389 168 0 1 64
0 5
0
0 0 20736 90
9 Direct In
-73 -6 -10 2
2 T2
-49 -16 -35 -8
0
0
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
1 T
6423 0 0
0
0
7 Ground~
168 412 289 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
3623 0 0
0
0
7 Ground~
168 297 236 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
8523 0 0
0
0
7 Ground~
168 199 347 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
3 GND
9623 0 0
0
0
2 +V
167 193 261 0 1 64
0 112
0
0 0 53600 46260
4 -15V
-13 2 15 10
3 V15
-10 -8 11 0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
9468 0 0
0
0
2 +V
167 193 177 0 1 64
0 113
0
0 0 53600 0
4 +15V
-13 -15 15 -7
3 V16
-10 -25 11 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
9254 0 0
0
0
8 Op-Amp5~
219 193 215 0 5 64
0 110 108 113 112 109
8 Op-Amp5~
0 0 17216 0
5 LF357
10 -13 45 -5
3 IC1
17 -23 38 -15
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 -33686019
88 -1 258 0 1 0 0 0
1 U
5587 0 0
0
0
12 TwistedPair~
219 64 215 0 4 64
0 124 125 115 114
12 TwistedPair~
0 0 16640 0
12 Twisted Pair
-41 -18 43 -10
5 CABL3
-17 -28 18 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -33686019
0 0 254 512 1 0 0 0
4 CABL
3333 0 0
0
0
5 Coax~
219 350 219 0 4 64
0 111 2 5 126
5 Coax~
0 0 16640 0
12 Coax Cable 2
-42 -20 42 -12
5 CABL4
-18 -30 17 -22
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 -33686019
0 0 252 512 1 0 0 0
4 CABL
619 0 0
0
0
10 Capacitor~
219 228 303 0 2 64
0 2 110
10 Capacitor~
0 0 17216 90
4 82pF
12 0 40 8
3 C24
15 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
4641 0 0
0
0
10 Capacitor~
219 207 107 0 2 64
0 108 109
10 Capacitor~
0 0 17216 0
4 82pF
-14 -18 14 -10
3 C23
-11 -28 10 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
5734 0 0
0
0
13 Var Resistor~
219 416 259 0 3 64
0 5 107 2
13 Var Resistor~
0 0 17216 23685390
7 10k 40%
-52 -5 -3 3
3 R43
-38 -15 -17 -7
0
0
30 %DA %1 %2 4000
%DB %2 %3 6000
0
0
4 SIP3
7

0 1 2 3 1 2 3 -33686019
82 0 272 0 1 0 0 0
1 R
3505 0 0
0
0
10 Capacitor~
219 499 259 0 2 64
0 2 103
10 Capacitor~
0 0 832 0
5 .01uF
-18 -18 17 -10
3 C21
-11 -28 10 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
7357 0 0
0
0
10 Capacitor~
219 507 115 0 2 64
0 101 7
10 Capacitor~
0 0 832 0
4 82pF
-14 -18 14 -10
3 C20
-11 -28 10 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
5588 0 0
0
0
12 NPN Trans:C~
219 664 248 0 3 64
0 89 96 100
12 NPN Trans:C~
0 0 832 0
6 MPSA06
18 0 60 8
2 Q3
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
81 -1 261 0 1 0 0 0
1 Q
3512 0 0
0
0
12 PNP Trans:C~
219 662 513 0 3 64
0 87 96 93
12 PNP Trans:C~
0 0 832 46772
6 MPSA56
18 0 60 8
2 Q4
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
113 0 262 0 1 0 0 0
1 Q
6225 0 0
0
0
12 PNP Trans:C~
219 794 515 0 3 64
0 90 48 92
12 PNP Trans:C~
0 0 832 46260
6 MPSA56
-64 0 -22 8
2 Q7
-50 -10 -36 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
113 0 262 0 1 0 0 0
1 Q
4624 0 0
0
0
11 Regulator3~
219 716 325 0 3 64
0 98 97 59
11 Regulator3~
0 0 832 23685390
5 LM334
-15 -8 20 0
3 IC3
-8 -17 13 -9
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
88 0 238 0 1 1 0 0
1 U
7815 0 0
0
0
10 Capacitor~
219 615 165 0 2 64
0 2 83
10 Capacitor~
0 0 832 90
5 100uF
11 0 46 8
2 C4
22 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
3296 0 0
0
0
12 N-EMOS 3T:A~
219 946 343 0 3 64
0 73 84 67
12 N-EMOS 3T:A~
0 0 832 512
6 IRF510
-6 -26 36 -18
3 Q24
4 -36 25 -28
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-220
7

0 2 1 3 2 1 3 -33686019
77 0 546 256 1 0 0 0
1 Q
6818 0 0
0
0
10 Capacitor~
219 881 341 0 2 64
0 67 73
10 Capacitor~
0 0 832 90
4 .1uF
12 0 40 8
2 C5
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
3184 0 0
0
0
13 Var Resistor~
219 990 282 0 3 64
0 73 73 84
13 Var Resistor~
0 0 832 23685390
7 10k 40%
-50 -4 -1 4
3 R18
-36 -15 -15 -7
0
0
30 %DA %1 %2 4000
%DB %2 %3 6000
0
0
4 SIP3
7

0 1 2 3 1 2 3 -33686019
82 0 272 0 1 0 0 0
1 R
7645 0 0
0
0
10 Capacitor~
219 877 271 0 2 64
0 2 85
10 Capacitor~
0 0 832 90
6 1500pF
12 0 54 8
3 C18
22 -10 43 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
8304 0 0
0
0
11 Regulator3~
219 1052 51 0 3 64
0 83 82 81
11 Regulator3~
0 0 4928 0
6 LM317T
-21 -28 21 -20
3 IC8
-11 -38 10 -30
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-220
7

0 3 1 2 3 1 2 -33686019
88 0 238 0 1 0 0 0
1 U
9203 0 0
0
0
10 Capacitor~
219 1169 743 0 2 64
0 60 54
10 Capacitor~
0 0 832 0
3 1uF
-11 -18 10 -10
3 C19
-11 -28 10 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
3686 0 0
0
0
8 Op-Amp5~
219 1321 737 0 5 64
0 54 53 52 2 55
8 Op-Amp5~
0 0 832 0
5 LM339
10 -14 45 -6
3 IC4
16 -24 37 -16
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 -33686019
88 -1 258 0 1 0 0 0
2 IC
3197 0 0
0
0
8 Caution~
219 1099 576 0 1 64
0 0
8 Caution~
0 0 49248 0
0
0
0
0
0
0
0
0
3

0 0 0 -33686019
0 0 721 0 1 0 0 0
3 SYM
7910 0 0
0
0
12 Zener Diode~
219 1469 599 0 2 64
0 26 38
12 Zener Diode~
0 0 832 90
7 1N4742A
13 1 62 9
2 D5
31 -10 45 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
100 0 281 0 1 0 0 0
1 D
5522 0 0
0
0
12 N-EMOS 3T:A~
219 1581 596 0 3 64
0 25 50 26
12 N-EMOS 3T:A~
0 0 832 0
7 IRFP240
-25 42 24 50
3 Q20
-11 31 10 39
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
77 0 546 0 1 0 0 0
1 Q
3636 0 0
0
0
10 Capacitor~
219 1451 420 0 2 64
0 48 29
10 Capacitor~
0 0 832 0
4 82pF
-14 -18 14 -10
2 C7
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
975 0 0
0
0
10 Capacitor~
219 1446 274 0 2 64
0 49 29
10 Capacitor~
0 0 832 0
5 150pF
-18 -18 17 -10
2 C6
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
7668 0 0
0
0
8 Op-Amp5~
219 1494 444 0 5 64
0 43 45 46 47 44
8 Op-Amp5~
0 0 832 180
5 LF411
-40 14 -5 22
3 IC5
-34 4 -13 12
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 8 4 6 3 2 8 4
6 -33686019
88 -1 258 0 1 0 0 0
1 U
3890 0 0
0
0
10 Capacitor~
219 1410 478 0 2 64
0 44 45
10 Capacitor~
0 0 832 0
5 .22uF
-18 -18 17 -10
2 C8
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
3461 0 0
0
0
10 Capacitor~
219 1575 438 0 2 64
0 43 2
10 Capacitor~
0 0 832 0
5 .22uF
-18 -18 17 -10
2 C9
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
8162 0 0
0
0
12 P-EMOS 3T:A~
219 1581 87 0 3 64
0 25 42 33
12 P-EMOS 3T:A~
0 0 832 46772
8 IRFP9240
-63 -24 -7 -16
3 Q16
-45 -34 -24 -26
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
109 0 552 0 1 0 0 0
1 Q
4417 0 0
0
0
6 Diode~
219 1727 378 0 2 64
0 31 32
6 Diode~
0 0 832 90
6 1N4002
12 0 54 8
3 D14
22 -10 43 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 -1 280 0 1 0 0 0
1 D
330 0 0
0
0
12 N-EMOS 3T:A~
219 1793 427 0 3 64
0 31 20 2
12 N-EMOS 3T:A~
0 0 832 0
8 VN0610LL
18 0 74 8
3 Q25
35 -10 56 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
77 0 546 0 1 0 0 0
1 Q
9669 0 0
0
0
12 Zener Diode~
219 1729 468 0 2 64
0 2 20
12 Zener Diode~
0 0 832 90
7 1N4742A
13 -2 62 6
3 D15
27 -12 48 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
100 0 281 0 1 0 0 0
1 D
5704 0 0
0
0
10 Capacitor~
219 1675 490 0 2 64
0 20 2
10 Capacitor~
0 0 832 0
4 10uF
-14 -18 14 -10
3 C10
-11 -28 10 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
3504 0 0
0
0
5 Fuse~
219 1994 42 0 2 64
0 33 28
5 Fuse~
0 0 4928 0
3 10A
-10 -16 11 -8
2 F1
-7 -26 7 -18
0
0
11 %D %1 %2 %S
0
0
4 FUSE
5

0 1 2 1 2 -33686019
88 0 246 0 1 0 0 0
1 F
3413 0 0
0
0
10 Capacitor~
219 1966 651 0 2 64
0 2 26
10 Capacitor~
0 0 832 90
4 .1uF
12 0 40 8
3 C14
15 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
9722 0 0
0
0
10 Capacitor~
219 2028 651 0 2 64
0 2 26
10 Capacitor~
0 0 832 90
5 100uF
11 0 46 8
3 C15
18 -10 39 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -33686019
67 -1 273 0 1 0 0 0
1 C
9512 0 0
0
0
12 Zener Diode~
219 1998 166 0 2 64
0 19 14
12 Zener Diode~
0 0 832 90
7 1N4742A
13 -2 62 6
3 D11
27 -12 48 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
100 0 281 0 1 0 0 0
1 D
7895 0 0
0
0
12 Zener Diode~
219 1998 222 0 2 64
0 19 2
12 Zener Diode~
0 0 832 23685390
7 1N4742A
13 -2 62 6
3 D10
27 -12 48 -4
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
100 0 281 0 1 0 0 0
1 D
6702 0 0
0
0
10 Polar Cap~
219 2069 156 0 2 64
0 14 2
10 Polar Cap~
0 0 832 23685390
4 10uF
11 4 39 12
3 C11
14 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 -1 274 0 1 0 0 0
1 C
3798 0 0
0
0
9 Resistor~
219 738 33 0 64 64
0 9 8 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
9 Resistor~
0 0 17248 0
5 5.11k
-17 -14 18 -6
3 R78
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 -1 271 0 1 0 0 0
1 R
3439 0 0
0
0
9 Resistor~
219 2233 229 0 2 64
0 24 23
9 Resistor~
0 0 864 0
2 1k
-7 -14 7 -6
3 R49
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
8595 0 0
0
0
9 Resistor~
219 2233 132 0 2 64
0 22 21
9 Resistor~
0 0 864 0
2 1k
-7 -14 7 -6
3 R50
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9295 0 0
0
0
9 Resistor~
219 1894 163 0 2 64
0 34 35
9 Resistor~
0 0 864 90
3 200
7 0 28 8
3 R64
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
8457 0 0
0
0
9 Resistor~
219 1775 163 0 2 64
0 34 36
9 Resistor~
0 0 864 90
3 200
7 0 28 8
3 R63
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
7780 0 0
0
0
9 Resistor~
219 1655 163 0 2 64
0 34 37
9 Resistor~
0 0 864 90
3 200
7 0 28 8
3 R62
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
5962 0 0
0
0
9 Resistor~
219 1894 579 0 2 64
0 39 38
9 Resistor~
0 0 864 90
3 200
7 0 28 8
3 R68
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3156 0 0
0
0
9 Resistor~
219 1775 579 0 2 64
0 40 38
9 Resistor~
0 0 864 90
3 200
7 0 28 8
3 R67
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9206 0 0
0
0
9 Resistor~
219 1655 579 0 2 64
0 41 38
9 Resistor~
0 0 864 90
3 200
7 0 28 8
3 R66
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
6360 0 0
0
0
9 Resistor~
219 1281 698 0 4 64
0 53 52 0 1
9 Resistor~
0 0 864 90
3 15k
7 0 28 8
3 R58
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3720 0 0
0
0
9 Resistor~
219 1334 415 0 2 64
0 63 49
9 Resistor~
0 0 864 90
2 1k
11 0 25 8
3 R31
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
6565 0 0
0
0
9 Resistor~
219 1040 413 0 4 64
0 65 2 0 -1
9 Resistor~
0 0 864 90
2 1k
11 0 25 8
3 R21
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
6565 0 0
0
0
9 Resistor~
219 1334 72 0 2 64
0 71 33
9 Resistor~
0 0 864 90
2 1k
11 0 25 8
3 R29
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
8521 0 0
0
0
9 Resistor~
219 1402 153 0 3 64
0 2 69 -1
9 Resistor~
0 0 864 90
2 2k
11 0 25 8
3 R33
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
578 0 0
0
0
9 Resistor~
219 1111 273 0 4 64
0 77 75 0 1
9 Resistor~
0 0 864 90
5 5.11k
7 0 42 8
3 R22
14 -10 35 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3756 0 0
0
0
9 Resistor~
219 1034 336 0 3 64
0 2 78 -1
9 Resistor~
0 0 864 90
2 1k
11 0 25 8
3 R20
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3435 0 0
0
0
9 Resistor~
219 1216 295 0 2 64
0 76 72
9 Resistor~
0 0 864 0
2 1k
-7 -14 7 -6
3 R23
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
822 0 0
0
0
9 Resistor~
219 1193 320 0 3 64
0 74 76 1
9 Resistor~
0 0 864 90
3 20k
7 0 28 8
3 R24
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3541 0 0
0
0
9 Resistor~
219 1220 359 0 3 64
0 74 66 1
9 Resistor~
0 0 864 0
3 10k
-10 -14 11 -6
3 R55
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
5454 0 0
0
0
9 Resistor~
219 1106 42 0 2 64
0 81 33
9 Resistor~
0 0 864 0
3 330
-10 -14 11 -6
3 R25
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
4961 0 0
0
0
9 Resistor~
219 1108 99 0 4 64
0 82 2 0 -1
9 Resistor~
0 0 864 0
5 27.4k
-17 -14 18 -6
3 R70
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
5218 0 0
0
0
9 Resistor~
219 785 587 0 3 64
0 59 90 1
9 Resistor~
0 0 864 90
3 10k
-26 0 -5 8
3 R10
-26 -10 -5 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
4436 0 0
0
0
9 Resistor~
219 679 586 0 3 64
0 59 87 1
9 Resistor~
0 0 864 90
3 10k
7 0 28 8
2 R1
10 -10 24 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9121 0 0
0
0
9 Resistor~
219 786 168 0 4 64
0 91 83 0 1
9 Resistor~
0 0 864 90
3 10k
-27 -1 -6 7
2 R7
-23 -11 -9 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9298 0 0
0
0
9 Resistor~
219 694 482 0 2 64
0 93 94
9 Resistor~
0 0 864 0
3 100
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9759 0 0
0
0
9 Resistor~
219 759 482 0 2 64
0 94 92
9 Resistor~
0 0 864 0
3 100
-10 -14 11 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
7712 0 0
0
0
9 Resistor~
219 677 412 0 2 64
0 94 95
9 Resistor~
0 0 864 0
5 33.2k
-17 -14 18 -6
3 R13
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
6691 0 0
0
0
9 Resistor~
219 761 288 0 2 64
0 98 99
9 Resistor~
0 0 864 0
3 100
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9275 0 0
0
0
9 Resistor~
219 598 374 0 2 64
0 105 96
9 Resistor~
0 0 864 0
5 2.05k
-17 -14 18 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3379 0 0
0
0
9 Resistor~
219 460 319 0 2 64
0 104 101
9 Resistor~
0 0 864 90
5 46.4k
7 0 42 8
3 R73
14 -10 35 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
373 0 0
0
0
9 Resistor~
219 540 374 0 2 64
0 106 105
9 Resistor~
0 0 864 0
5 2.05k
-17 -14 18 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
4818 0 0
0
0
9 Resistor~
219 508 401 0 3 64
0 2 106 -1
9 Resistor~
0 0 864 90
5 46.4k
7 0 42 8
2 R8
18 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
6965 0 0
0
0
9 Resistor~
219 144 209 0 2 64
0 115 108
9 Resistor~
0 0 17248 0
5 46.4k
-17 -14 18 -6
3 R75
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3783 0 0
0
0
9 Resistor~
219 144 221 0 2 64
0 114 110
9 Resistor~
0 0 17248 0
5 46.4k
-18 18 17 26
3 R76
-11 7 10 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
8577 0 0
0
0
9 Resistor~
219 168 305 0 3 64
0 2 110 -1
9 Resistor~
0 0 17248 90
5 46.4k
7 0 42 8
3 R41
14 -10 35 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
410 0 0
0
0
9 Resistor~
219 271 215 0 2 64
0 109 111
9 Resistor~
0 0 17248 0
3 402
-10 -14 11 -6
3 R42
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
5148 0 0
0
0
9 Resistor~
219 205 148 0 2 64
0 108 109
9 Resistor~
0 0 17248 0
5 46.4k
-17 -14 18 -6
3 R77
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
4242 0 0
0
0
9 Resistor~
219 506 77 0 2 64
0 101 7
9 Resistor~
0 0 864 0
5 46.4k
-17 -14 18 -6
3 R74
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3163 0 0
0
0
9 Resistor~
219 695 288 0 2 64
0 100 98
9 Resistor~
0 0 864 0
3 100
-10 -14 11 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3470 0 0
0
0
9 Resistor~
219 673 328 0 3 64
0 59 97 1
9 Resistor~
0 0 864 0
5 33.2k
-17 -14 18 -6
3 R12
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
5476 0 0
0
0
9 Resistor~
219 669 166 0 4 64
0 89 83 0 1
9 Resistor~
0 0 864 90
3 10k
7 0 28 8
3 R11
8 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3680 0 0
0
0
9 Resistor~
219 936 166 0 4 64
0 88 83 0 1
9 Resistor~
0 0 864 90
2 1k
11 0 25 8
3 R15
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
4465 0 0
0
0
9 Resistor~
219 936 586 0 3 64
0 59 86 1
9 Resistor~
0 0 864 90
2 1k
11 0 25 8
3 R16
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
344 0 0
0
0
9 Resistor~
219 906 246 0 2 64
0 85 73
9 Resistor~
0 0 864 0
3 402
-10 -14 11 -6
3 R17
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3539 0 0
0
0
9 Resistor~
219 986 436 0 2 64
0 67 84
9 Resistor~
0 0 864 90
5 5.11k
7 0 42 8
3 R19
14 -10 35 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3669 0 0
0
0
9 Resistor~
219 1053 137 0 3 64
0 83 80 1
9 Resistor~
0 0 864 0
3 100
-10 -14 11 -6
3 R26
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3321 0 0
0
0
9 Resistor~
219 1013 99 0 3 64
0 83 82 1
9 Resistor~
0 0 864 0
5 1.21k
-17 -14 18 -6
3 R69
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
350 0 0
0
0
9 Resistor~
219 1334 291 0 2 64
0 49 64
9 Resistor~
0 0 864 90
2 1k
11 0 25 8
3 R30
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
932 0 0
0
0
9 Resistor~
219 1268 589 0 2 64
0 54 66
9 Resistor~
0 0 864 90
2 1k
11 0 25 8
3 R56
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
5914 0 0
0
0
9 Resistor~
219 1174 557 0 3 64
0 59 61 1
9 Resistor~
0 0 864 0
3 100
-10 -14 11 -6
3 R28
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
4398 0 0
0
0
9 Resistor~
219 1060 677 0 3 64
0 59 58 1
9 Resistor~
0 0 864 0
5 1.12k
-17 -14 18 -6
3 R71
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
6628 0 0
0
0
9 Resistor~
219 1100 711 0 2 64
0 60 58
9 Resistor~
0 0 864 90
5 27.4k
7 0 42 8
3 R72
14 -10 35 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9418 0 0
0
0
9 Resistor~
219 1173 620 0 2 64
0 57 26
9 Resistor~
0 0 864 0
3 330
-10 -14 11 -6
3 R27
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9849 0 0
0
0
9 Resistor~
219 1334 599 0 2 64
0 26 51
9 Resistor~
0 0 864 90
2 1k
11 0 25 8
3 R32
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
4899 0 0
0
0
9 Resistor~
219 1218 697 0 4 64
0 54 52 0 1
9 Resistor~
0 0 864 90
4 825k
8 0 36 8
3 R57
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3179 0 0
0
0
9 Resistor~
219 1380 713 0 2 64
0 55 56
9 Resistor~
0 0 864 90
5 2.05k
7 0 42 8
3 R60
14 -10 35 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
898 0 0
0
0
9 Resistor~
219 1281 776 0 3 64
0 2 53 -1
9 Resistor~
0 0 864 90
3 15k
7 0 28 8
3 R59
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 1402 533 0 4 64
0 38 2 0 -1
9 Resistor~
0 0 864 90
2 2k
11 0 25 8
3 R34
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
4185 0 0
0
0
9 Resistor~
219 1536 579 0 2 64
0 50 38
9 Resistor~
0 0 864 90
3 200
7 0 28 8
3 R65
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
8302 0 0
0
0
9 Resistor~
219 1449 381 0 2 64
0 48 29
9 Resistor~
0 0 864 0
5 5.11k
-17 -14 18 -6
3 R37
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9670 0 0
0
0
9 Resistor~
219 1447 313 0 2 64
0 49 29
9 Resistor~
0 0 864 0
4 1.5k
-14 -14 14 -6
3 R36
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3998 0 0
0
0
9 Resistor~
219 1353 338 0 3 64
0 2 49 -1
9 Resistor~
0 0 864 90
2 50
11 0 25 8
3 R35
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
7488 0 0
0
0
9 Resistor~
219 1378 408 0 2 64
0 44 48
9 Resistor~
0 0 864 90
3 10k
7 0 28 8
3 R38
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9634 0 0
0
0
9 Resistor~
219 1555 478 0 4 64
0 45 2 0 -1
9 Resistor~
0 0 864 0
4 825k
-14 -14 14 -6
3 R40
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
6103 0 0
0
0
9 Resistor~
219 1521 411 0 2 64
0 43 29
9 Resistor~
0 0 864 90
4 825k
8 0 36 8
3 R39
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
9627 0 0
0
0
9 Resistor~
219 1536 163 0 2 64
0 34 42
9 Resistor~
0 0 864 90
3 200
7 0 28 8
3 R61
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
5925 0 0
0
0
9 Resistor~
219 1673 396 0 4 64
0 20 32 0 1
9 Resistor~
0 0 864 90
4 825k
8 0 36 8
3 R51
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
82 0 0
0
0
9 Resistor~
219 1905 431 0 3 64
0 2 30 -1
9 Resistor~
0 0 864 90
2 1k
11 0 25 8
3 R52
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3195 0 0
0
0
9 Resistor~
219 1973 138 0 2 64
0 25 14
9 Resistor~
0 0 864 0
4 825k
-14 -14 14 -6
3 R44
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
8459 0 0
0
0
9 Resistor~
219 2120 168 0 3 64
0 2 18 -1
9 Resistor~
0 0 864 90
2 1k
11 0 25 8
3 R45
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
3620 0 0
0
0
9 Resistor~
219 2120 99 0 4 64
0 18 17 0 1
9 Resistor~
0 0 864 90
5 5.11k
7 0 42 8
3 R46
14 -10 35 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
344 0 0
0
0
9 Resistor~
219 2168 273 0 4 64
0 15 13 0 1
9 Resistor~
0 0 864 0
5 5.11k
-17 -14 18 -6
3 R48
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
6142 0 0
0
0
9 Resistor~
219 2107 273 0 3 64
0 2 15 -1
9 Resistor~
0 0 864 0
2 1k
-7 -14 7 -6
3 R47
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 0 0 0
1 R
6317 0 0
0
0
279
0 0 6 0 0 4480 0 0 0 0 0 5
583 3
895 3
895 120
583 120
583 3
2 1 7 0 0 4096 0 172 7 0 0 4
524 77
643 77
643 78
655 78
2 2 8 0 0 4224 0 135 4 0 0 2
756 33
774 33
2 1 9 0 0 4224 0 1 135 0 0 2
698 33
720 33
1 1 2 0 0 4096 0 1 79 0 0 3
678 33
641 33
641 49
1 1 10 0 0 4224 0 4 2 0 0 3
808 37
829 37
829 31
3 2 11 0 0 8320 0 7 5 0 0 4
751 78
761 78
761 49
774 49
1 1 3 0 0 4224 0 3 5 0 0 2
816 53
808 53
2 1 2 0 0 0 0 7 6 0 0 3
655 86
649 86
649 97
0 0 12 0 0 12672 0 0 0 0 0 5
16 71
448 71
448 409
14 409
14 71
2 1 13 0 0 4224 0 206 8 0 0 2
2186 273
2198 273
2 0 14 0 0 8192 0 16 0 0 26 3
2148 223
2112 223
2112 138
1 0 15 0 0 8320 0 16 0 0 14 3
2148 235
2136 235
2136 273
2 1 15 0 0 0 0 207 206 0 0 2
2125 273
2150 273
1 0 2 0 0 4096 0 207 0 0 23 2
2089 273
1998 273
1 3 16 0 0 4224 0 9 15 0 0 2
2166 88
2166 119
1 2 17 0 0 4224 0 10 205 0 0 2
2120 73
2120 81
1 0 2 0 0 0 0 204 0 0 21 3
2120 186
2120 198
2068 198
2 0 18 0 0 4096 0 15 0 0 20 2
2148 126
2120 126
1 2 18 0 0 4224 0 205 204 0 0 2
2120 117
2120 150
2 0 2 0 0 4096 0 134 0 0 15 2
2068 163
2068 273
1 0 14 0 0 0 0 134 0 0 26 2
2068 146
2068 138
2 1 2 0 0 0 0 133 11 0 0 2
1998 232
1998 282
1 1 19 0 0 4224 0 132 133 0 0 2
1998 176
1998 212
2 0 14 0 0 0 0 132 0 0 26 2
1998 156
1998 138
2 1 14 0 0 4224 0 203 15 0 0 2
1991 138
2148 138
1 1 2 0 0 0 0 12 13 0 0 4
2262 66
2262 59
2315 59
2315 68
1 0 20 0 0 4096 0 17 0 0 34 2
2289 132
2315 132
2 2 21 0 0 4224 0 137 17 0 0 2
2251 132
2269 132
5 1 22 0 0 4224 0 15 137 0 0 2
2184 132
2215 132
1 0 20 0 0 0 0 14 0 0 34 2
2290 229
2315 229
2 2 23 0 0 4224 0 136 14 0 0 2
2251 229
2270 229
5 1 24 0 0 4224 0 16 136 0 0 2
2184 229
2215 229
1 2 20 0 0 12416 0 128 13 0 0 5
1666 490
1646 490
1646 301
2315 301
2315 102
1 0 25 0 0 4096 0 203 0 0 64 2
1955 138
1945 138
1 1 2 0 0 0 0 19 130 0 0 2
1966 675
1966 660
1 1 2 0 0 0 0 18 131 0 0 2
2028 675
2028 660
2 0 26 0 0 4096 0 131 0 0 128 2
2028 642
2028 620
2 0 26 0 0 0 0 130 0 0 128 2
1966 642
1966 620
2 1 27 0 0 4224 0 21 20 0 0 2
2093 620
2106 620
2 1 28 0 0 4224 0 129 22 0 0 2
2016 42
2029 42
3 1 4 0 0 4224 0 28 23 0 0 2
1849 351
1961 351
0 1 29 0 0 4224 0 0 28 100 0 4
1521 313
1868 313
1868 344
1849 344
1 1 2 0 0 0 0 202 24 0 0 2
1905 449
1905 464
2 2 30 0 0 4224 0 25 202 0 0 3
1884 398
1905 398
1905 413
1 0 31 0 0 4096 0 25 0 0 57 2
1864 398
1799 398
1 0 31 0 0 8320 0 125 0 0 57 3
1727 388
1727 398
1799 398
1 0 32 0 0 4096 0 27 0 0 56 2
1780 347
1780 357
2 0 20 0 0 0 0 127 0 0 51 2
1729 458
1729 436
1 0 20 0 0 0 0 201 0 0 51 2
1673 414
1673 436
2 0 20 0 0 0 0 126 0 0 34 2
1775 436
1646 436
1 0 2 0 0 0 0 127 0 0 53 2
1729 478
1729 490
2 0 2 0 0 4224 0 128 0 0 54 2
1684 490
1799 490
3 1 2 0 0 0 0 126 26 0 0 2
1799 445
1799 507
2 0 32 0 0 4096 0 125 0 0 56 2
1727 368
1727 357
2 4 32 0 0 8320 0 201 28 0 0 3
1673 378
1673 357
1819 357
5 1 31 0 0 0 0 28 126 0 0 3
1819 381
1799 381
1799 409
1 0 25 0 0 4096 0 33 0 0 60 2
1826 578
1826 537
1 0 25 0 0 4096 0 34 0 0 60 2
1706 579
1706 537
1 0 25 0 0 8192 0 118 0 0 64 3
1587 578
1587 537
1945 537
1 0 25 0 0 0 0 30 0 0 63 2
1826 105
1826 199
1 0 25 0 0 0 0 31 0 0 63 2
1706 105
1706 199
1 0 25 0 0 0 0 124 0 0 64 3
1587 105
1587 199
1945 199
1 1 25 0 0 4224 0 29 32 0 0 2
1945 105
1945 578
3 0 33 0 0 4096 0 29 0 0 181 2
1945 69
1945 42
3 0 33 0 0 0 0 30 0 0 181 2
1826 69
1826 42
3 0 33 0 0 0 0 31 0 0 181 2
1706 69
1706 42
1 0 34 0 0 4096 0 140 0 0 84 2
1655 181
1655 224
1 0 34 0 0 0 0 139 0 0 84 2
1775 181
1775 224
2 2 35 0 0 4224 0 138 29 0 0 3
1894 145
1894 78
1921 78
2 2 36 0 0 4224 0 139 30 0 0 3
1775 145
1775 78
1802 78
2 2 37 0 0 4224 0 140 31 0 0 3
1655 145
1655 78
1682 78
2 0 38 0 0 4096 0 142 0 0 111 2
1775 561
1775 555
2 0 38 0 0 0 0 143 0 0 111 2
1655 561
1655 555
3 0 26 0 0 0 0 34 0 0 128 2
1706 615
1706 620
3 0 26 0 0 0 0 33 0 0 128 2
1826 614
1826 620
3 0 26 0 0 0 0 32 0 0 128 2
1945 614
1945 620
1 2 39 0 0 8320 0 141 32 0 0 3
1894 597
1894 605
1921 605
1 2 40 0 0 8320 0 142 33 0 0 3
1775 597
1775 605
1802 605
1 2 41 0 0 8320 0 143 34 0 0 3
1655 597
1655 606
1682 606
1 0 34 0 0 0 0 200 0 0 84 2
1536 181
1536 224
3 0 33 0 0 0 0 124 0 0 181 2
1587 69
1587 42
2 2 42 0 0 4224 0 200 124 0 0 3
1536 145
1536 78
1563 78
1 1 34 0 0 8320 0 35 138 0 0 4
1469 141
1469 224
1894 224
1894 181
2 0 33 0 0 4096 0 35 0 0 181 2
1469 121
1469 42
2 0 2 0 0 0 0 198 0 0 87 2
1573 478
1590 478
2 1 2 0 0 0 0 123 36 0 0 3
1584 438
1590 438
1590 487
1 0 43 0 0 4096 0 199 0 0 89 2
1521 429
1521 438
1 1 43 0 0 4224 0 121 123 0 0 2
1512 438
1566 438
1 0 44 0 0 8192 0 122 0 0 95 3
1401 478
1378 478
1378 444
2 0 45 0 0 8192 0 121 0 0 92 3
1512 450
1521 450
1521 478
2 1 45 0 0 4224 0 122 198 0 0 2
1419 478
1537 478
1 3 46 0 0 4224 0 37 121 0 0 2
1494 487
1494 457
1 4 47 0 0 4224 0 38 121 0 0 2
1494 423
1494 431
5 1 44 0 0 4224 0 121 197 0 0 3
1476 444
1378 444
1378 426
2 0 29 0 0 0 0 119 0 0 105 3
1460 420
1475 420
1475 381
1 0 48 0 0 8192 0 119 0 0 191 3
1442 420
1422 420
1422 381
2 0 48 0 0 0 0 197 0 0 191 2
1378 390
1378 381
2 0 29 0 0 0 0 120 0 0 100 3
1455 274
1475 274
1475 313
2 2 29 0 0 0 0 195 199 0 0 3
1465 313
1521 313
1521 393
1 1 2 0 0 0 0 196 39 0 0 2
1353 356
1353 362
2 0 49 0 0 4096 0 196 0 0 103 2
1353 320
1353 313
0 0 49 0 0 4096 0 0 0 141 104 2
1334 313
1421 313
1 1 49 0 0 0 0 120 195 0 0 4
1437 274
1421 274
1421 313
1429 313
2 0 29 0 0 0 0 194 0 0 100 2
1467 381
1521 381
3 0 26 0 0 0 0 118 0 0 128 2
1587 614
1587 620
1 2 50 0 0 8320 0 193 118 0 0 3
1536 597
1536 605
1563 605
2 0 38 0 0 0 0 193 0 0 111 2
1536 561
1536 555
1 0 26 0 0 0 0 117 0 0 128 2
1469 609
1469 620
2 0 38 0 0 4096 0 117 0 0 111 2
1469 589
1469 555
0 2 38 0 0 4224 0 0 141 112 0 3
1402 555
1894 555
1894 561
1 3 38 0 0 0 0 192 41 0 0 2
1402 551
1402 560
2 1 2 0 0 0 0 192 40 0 0 4
1402 515
1402 513
1452 513
1452 517
1 0 26 0 0 4096 0 41 0 0 128 2
1402 596
1402 620
0 2 51 0 0 4224 0 0 41 129 0 2
1334 578
1379 578
1 0 52 0 0 8192 0 42 0 0 124 3
1380 670
1380 665
1321 665
1 0 2 0 0 0 0 191 0 0 121 3
1281 794
1281 800
1321 800
2 0 53 0 0 4096 0 115 0 0 119 2
1303 731
1281 731
1 2 53 0 0 4224 0 144 191 0 0 2
1281 716
1281 758
2 0 52 0 0 0 0 144 0 0 122 2
1281 680
1281 665
4 1 2 0 0 0 0 115 44 0 0 2
1321 750
1321 806
2 0 52 0 0 8320 0 189 0 0 124 3
1218 679
1218 665
1321 665
1 0 54 0 0 4096 0 189 0 0 131 2
1218 715
1218 743
1 3 52 0 0 0 0 43 115 0 0 2
1321 657
1321 724
5 1 55 0 0 4224 0 115 190 0 0 3
1339 737
1380 737
1380 731
2 2 56 0 0 4224 0 42 190 0 0 2
1380 690
1380 695
1 0 26 0 0 0 0 188 0 0 128 2
1334 617
1334 620
2 1 26 0 0 4224 0 187 21 0 0 2
1191 620
2049 620
1 2 51 0 0 0 0 47 188 0 0 2
1334 575
1334 581
1 0 54 0 0 4224 0 183 0 0 131 2
1268 607
1268 743
2 1 54 0 0 0 0 114 115 0 0 2
1178 743
1303 743
3 1 57 0 0 4224 0 46 187 0 0 2
1128 620
1155 620
2 0 58 0 0 4096 0 185 0 0 136 2
1078 677
1100 677
1 0 59 0 0 8192 0 185 0 0 207 3
1042 677
1018 677
1018 620
1 1 60 0 0 8320 0 186 114 0 0 3
1100 729
1100 743
1160 743
2 2 58 0 0 4224 0 46 186 0 0 2
1100 653
1100 693
2 2 61 0 0 4224 0 184 47 0 0 2
1192 557
1311 557
1 0 59 0 0 4096 0 184 0 0 207 3
1156 557
1056 557
1056 620
1 3 62 0 0 4224 0 48 47 0 0 2
1334 530
1334 539
1 3 63 0 0 4224 0 145 48 0 0 2
1334 433
1334 494
1 2 49 0 0 4224 0 182 145 0 0 2
1334 309
1334 397
3 2 64 0 0 4224 0 55 182 0 0 2
1334 264
1334 273
2 0 65 0 0 4224 0 52 0 0 144 2
1088 436
1040 436
1 1 65 0 0 0 0 146 51 0 0 2
1040 431
1040 451
1 0 66 0 0 8192 0 52 0 0 151 3
1111 454
1111 466
1268 466
1 0 67 0 0 4096 0 50 0 0 190 2
1040 501
1040 512
3 0 2 0 0 0 0 52 0 0 149 2
1111 418
1111 392
2 2 68 0 0 4224 0 51 50 0 0 2
1040 471
1040 481
2 1 2 0 0 0 0 146 49 0 0 4
1040 395
1040 392
1132 392
1132 400
2 0 66 0 0 0 0 153 0 0 151 2
1238 359
1268 359
1 2 66 0 0 4224 0 58 183 0 0 2
1268 313
1268 571
3 1 2 0 0 0 0 58 53 0 0 4
1268 277
1268 257
1246 257
1246 263
1 0 33 0 0 0 0 56 0 0 181 2
1402 85
1402 42
2 0 33 0 0 0 0 147 0 0 181 2
1334 54
1334 42
3 2 69 0 0 4224 0 56 148 0 0 2
1402 121
1402 135
1 1 2 0 0 0 0 148 54 0 0 2
1402 171
1402 182
3 1 70 0 0 4224 0 57 55 0 0 2
1334 155
1334 228
2 0 71 0 0 4224 0 56 0 0 159 2
1379 103
1334 103
1 1 71 0 0 0 0 147 57 0 0 2
1334 90
1334 119
2 2 72 0 0 4224 0 151 58 0 0 2
1234 295
1245 295
2 0 73 0 0 4096 0 63 0 0 193 2
1034 257
1034 246
1 0 74 0 0 4224 0 152 0 0 163 2
1193 338
1193 359
1 1 74 0 0 0 0 59 153 0 0 2
1186 359
1202 359
1 2 75 0 0 4224 0 65 149 0 0 2
1111 236
1111 255
2 0 76 0 0 4096 0 152 0 0 166 2
1193 302
1193 295
2 1 76 0 0 4224 0 60 151 0 0 2
1186 295
1198 295
1 0 77 0 0 4224 0 60 0 0 168 2
1166 295
1111 295
1 3 77 0 0 0 0 149 62 0 0 2
1111 291
1111 300
2 0 78 0 0 4224 0 62 0 0 172 2
1088 318
1034 318
1 0 2 0 0 0 0 150 0 0 171 2
1034 354
1111 354
1 1 2 0 0 0 0 62 61 0 0 2
1111 336
1111 359
2 2 78 0 0 0 0 64 150 0 0 2
1034 304
1034 318
1 1 79 0 0 4224 0 63 64 0 0 2
1034 277
1034 284
2 2 80 0 0 4224 0 180 57 0 0 2
1071 137
1311 137
3 1 81 0 0 4224 0 113 154 0 0 2
1080 42
1088 42
2 0 33 0 0 0 0 67 0 0 181 2
1212 62
1212 42
2 0 33 0 0 0 0 68 0 0 181 2
1148 62
1148 42
1 0 2 0 0 0 0 68 0 0 179 2
1148 80
1148 99
2 0 2 0 0 0 0 155 0 0 180 2
1126 99
1212 99
1 1 2 0 0 0 0 67 66 0 0 2
1212 80
1212 107
2 1 33 0 0 4224 0 154 129 0 0 2
1124 42
1972 42
2 0 82 0 0 4096 0 113 0 0 183 2
1052 75
1052 99
2 1 82 0 0 4224 0 181 155 0 0 2
1031 99
1090 99
1 0 83 0 0 4096 0 181 0 0 185 2
995 99
984 99
1 0 83 0 0 8192 0 113 0 0 218 3
1024 42
984 42
984 137
2 0 84 0 0 4096 0 109 0 0 189 2
960 352
986 352
2 0 73 0 0 8192 0 111 0 0 193 3
998 276
1004 276
1004 246
1 0 67 0 0 4096 0 179 0 0 190 2
986 454
986 512
3 2 84 0 0 4224 0 111 179 0 0 2
986 296
986 418
0 2 67 0 0 4224 0 0 48 199 0 2
936 512
1311 512
0 1 48 0 0 4224 0 0 194 221 0 2
859 381
1431 381
1 0 73 0 0 0 0 111 0 0 193 2
986 260
986 246
0 2 73 0 0 4224 0 0 55 210 0 2
936 246
1311 246
2 0 73 0 0 0 0 178 0 0 210 2
924 246
936 246
1 1 2 0 0 0 0 112 69 0 0 2
877 280
877 290
1 2 85 0 0 8320 0 178 112 0 0 3
888 246
877 246
877 262
1 0 67 0 0 0 0 110 0 0 199 3
881 350
881 369
936 369
2 0 73 0 0 0 0 110 0 0 210 3
881 332
881 312
936 312
3 1 67 0 0 0 0 109 70 0 0 2
936 361
936 523
3 2 86 0 0 4224 0 70 177 0 0 2
936 559
936 568
1 0 59 0 0 0 0 177 0 0 207 2
936 604
936 620
2 0 87 0 0 4224 0 70 0 0 220 2
913 541
679 541
2 0 59 0 0 0 0 72 0 0 207 2
625 629
625 620
1 1 2 0 0 0 0 72 71 0 0 2
625 647
625 659
1 0 59 0 0 0 0 157 0 0 207 2
679 604
679 620
1 0 59 0 0 0 0 156 0 0 207 2
785 605
785 620
1 1 59 0 0 4224 0 73 46 0 0 2
609 620
1072 620
1 0 83 0 0 12288 0 77 0 0 218 4
728 384
728 376
849 376
849 137
0 0 59 0 0 0 0 0 0 233 207 3
738 364
839 364
839 620
1 1 73 0 0 0 0 74 109 0 0 2
936 229
936 325
2 0 83 0 0 0 0 176 0 0 218 2
936 148
936 137
3 1 88 0 0 4224 0 74 176 0 0 2
936 193
936 184
2 0 89 0 0 4224 0 74 0 0 222 2
913 211
669 211
1 1 2 0 0 0 0 108 75 0 0 2
615 174
615 187
2 0 83 0 0 0 0 108 0 0 218 2
615 156
615 137
2 0 83 0 0 0 0 175 0 0 218 2
669 148
669 137
2 0 83 0 0 0 0 158 0 0 218 2
786 150
786 137
1 1 83 0 0 4224 0 76 180 0 0 2
609 137
1035 137
1 2 90 0 0 4224 0 106 156 0 0 2
785 533
785 569
1 2 87 0 0 0 0 105 157 0 0 4
667 531
667 541
679 541
679 568
2 2 48 0 0 0 0 78 106 0 0 4
809 248
859 248
859 515
808 515
1 1 89 0 0 0 0 175 104 0 0 2
669 184
669 230
1 1 91 0 0 4224 0 158 78 0 0 2
786 186
786 230
2 3 92 0 0 8320 0 160 106 0 0 3
777 482
785 482
785 497
1 3 93 0 0 8320 0 159 105 0 0 3
676 482
667 482
667 495
0 0 94 0 0 4096 0 0 0 227 228 2
728 482
728 449
2 1 94 0 0 0 0 159 160 0 0 2
712 482
741 482
1 3 94 0 0 12416 0 161 77 0 0 5
659 412
651 412
651 449
728 449
728 440
2 2 95 0 0 4224 0 161 77 0 0 4
695 412
700 412
700 412
695 412
2 0 96 0 0 4096 0 163 0 0 231 2
616 374
634 374
2 2 96 0 0 8320 0 104 105 0 0 4
646 248
634 248
634 513
644 513
2 2 97 0 0 4224 0 174 107 0 0 4
691 328
700 328
700 328
695 328
1 3 59 0 0 0 0 174 107 0 0 7
655 328
651 328
651 364
738 364
738 364
728 364
728 356
1 0 98 0 0 4096 0 107 0 0 235 2
728 300
728 288
2 1 98 0 0 4224 0 173 162 0 0 2
713 288
743 288
3 2 99 0 0 4224 0 78 162 0 0 3
786 266
786 288
779 288
3 1 100 0 0 4224 0 104 173 0 0 3
669 266
669 288
677 288
1 0 101 0 0 4096 0 103 0 0 241 2
498 115
460 115
2 0 7 0 0 0 0 103 0 0 240 2
516 115
550 115
5 0 7 0 0 8320 0 83 0 0 2 3
537 208
550 208
550 77
1 0 101 0 0 8320 0 172 0 0 247 3
488 77
460 77
460 202
2 0 102 0 0 4096 0 80 0 0 249 2
507 180
519 180
1 0 2 0 0 0 0 80 0 0 246 3
489 180
477 180
477 214
2 0 103 0 0 4096 0 102 0 0 248 2
508 259
519 259
1 0 2 0 0 0 0 102 0 0 246 2
490 259
477 259
1 1 2 0 0 0 0 83 81 0 0 3
501 214
477 214
477 273
2 2 101 0 0 0 0 83 164 0 0 3
501 202
460 202
460 301
4 1 103 0 0 4224 0 83 84 0 0 2
519 221
519 272
1 3 102 0 0 4224 0 82 83 0 0 2
519 156
519 195
1 0 104 0 0 4096 0 164 0 0 251 2
460 337
460 374
3 1 104 0 0 8320 0 89 86 0 0 3
435 360
435 374
478 374
1 0 2 0 0 0 0 85 0 0 253 2
543 440
543 427
1 1 2 0 0 0 0 166 87 0 0 4
508 419
508 427
571 427
571 409
2 0 105 0 0 4096 0 87 0 0 256 2
571 391
571 374
2 0 106 0 0 4096 0 166 0 0 257 2
508 383
508 374
2 1 105 0 0 4224 0 165 163 0 0 2
558 374
580 374
2 1 106 0 0 4224 0 86 165 0 0 2
496 374
522 374
4 1 2 0 0 0 0 89 88 0 0 2
427 360
427 380
1 2 107 0 0 4224 0 89 101 0 0 3
435 264
435 253
424 253
3 0 5 0 0 4096 0 98 0 0 262 2
398 215
412 215
3 1 2 0 0 0 0 101 91 0 0 2
412 273
412 283
1 1 5 0 0 8320 0 90 101 0 0 3
400 166
412 166
412 237
1 0 108 0 0 4096 0 171 0 0 266 2
187 148
168 148
2 0 109 0 0 4096 0 171 0 0 265 2
223 148
242 148
2 0 109 0 0 8320 0 100 0 0 272 3
216 107
242 107
242 215
1 0 108 0 0 8320 0 100 0 0 276 3
198 107
168 107
168 209
2 1 2 0 0 0 0 98 92 0 0 3
302 223
297 223
297 230
1 0 2 0 0 0 0 93 0 0 269 2
199 341
199 327
1 1 2 0 0 0 0 169 99 0 0 4
168 323
168 327
228 327
228 312
2 0 110 0 0 8192 0 99 0 0 271 3
228 294
228 279
168 279
2 0 110 0 0 4224 0 169 0 0 277 2
168 287
168 221
5 1 109 0 0 0 0 96 170 0 0 2
211 215
253 215
2 1 111 0 0 4224 0 170 98 0 0 2
289 215
302 215
4 1 112 0 0 4224 0 96 94 0 0 2
193 228
193 246
1 3 113 0 0 4224 0 95 96 0 0 2
193 186
193 202
2 2 108 0 0 0 0 96 167 0 0 2
175 209
162 209
1 2 110 0 0 0 0 96 168 0 0 2
175 221
162 221
4 1 114 0 0 12416 0 97 168 0 0 4
112 219
118 219
118 221
126 221
3 1 115 0 0 12416 0 97 167 0 0 4
112 211
118 211
118 209
126 209
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 112
11 418 387 479
16 423 384 468
112 This schematic is configured so that items in 
Block A and Block B will not be included in the 
PCB netlist.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
584 0 645 23
589 5 642 20
7 Block B
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 32
662 84 788 121
666 88 785 116
32 Bridge output to 
next channel
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
14 69 75 92
19 74 72 89
7 Block A
-16 0 0 0 400 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 62
9 3 379 56
14 7 374 45
62 2 Channel Audio Amplifier
Schematic Only (not for simulation)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
864 804 1016 828
868 808 1012 824
18 Heat sink required
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
