CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 3
4 68 403 314
7 5.000 V
7 5.000 V
3 GND
4 68 403 314
42991616 0
0
0
0
0
0
0
7
14 Logic Display~
6 168 35 0 1 3
10 4
0
0 0 53296 0
6 100MEG
3 -16 45 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8953 0 0
0
0
7 Ground~
168 313 183 0 1 3
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
14 NO PushButton~
191 280 137 0 2 5
0 2 5
0
0 0 20576 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3618 0 0
0
0
14 NO PushButton~
191 209 128 0 2 5
0 2 6
0
0 0 20576 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
6153 0 0
0
0
8 Hex Key~
166 31 39 0 11 11
0 14 13 12 11 0 0 0 0 0
0 48
0
0 0 20512 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
5394 0 0
0
0
8 Hex Key~
166 71 39 0 11 11
0 10 9 8 7 0 0 0 0 0
3 51
0
0 0 20512 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7734 0 0
0
0
5 Delay
94 121 109 0 11 23
0 11 12 13 14 7 8 9 10 4
5 6
5 Delay
1 0 4224 0
0
0
0
0
0
0
0
0
23

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 0 0 0 0 0
0
9914 0 0
0
0
13
1 0 2 0 0 12416 0 4 0 0 2 4
226 136
242 136
242 159
313 159
1 1 2 0 0 0 0 3 2 0 0 3
297 145
313 145
313 177
1 9 4 0 0 4224 0 1 7 0 0 3
168 53
168 91
153 91
10 2 5 0 0 4224 0 7 3 0 0 2
159 145
263 145
11 2 6 0 0 4224 0 7 4 0 0 2
159 136
192 136
4 5 7 0 0 4224 0 6 7 0 0 3
62 63
62 118
89 118
3 6 8 0 0 4224 0 6 7 0 0 3
68 63
68 127
89 127
2 7 9 0 0 4224 0 6 7 0 0 3
74 63
74 136
89 136
1 8 10 0 0 4224 0 6 7 0 0 3
80 63
80 145
89 145
4 1 11 0 0 8320 0 5 7 0 0 3
22 63
22 82
89 82
3 2 12 0 0 8320 0 5 7 0 0 3
28 63
28 91
89 91
2 3 13 0 0 8320 0 5 7 0 0 3
34 63
34 100
89 100
1 4 14 0 0 8320 0 5 7 0 0 3
40 63
40 109
89 109
2
16 8 0 0 0 0 0 0 0 0 0 0 54
6 System
0 0 0 5
188 72 253 100
192 76 239 96
5 Reset
16 8 0 0 0 0 0 0 0 0 0 0 54
6 System
0 0 0 12
257 60 327 112
261 64 313 104
12 Start
Delay
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
