CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 800 319
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 800 319
9961490 0
0
6 Title:
5 Name:
0
0
0
7
7 Ground~
168 193 157 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
5 SAVE-
218 238 55 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
29 *Combine
*TRAN 0.000 10.00 0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
4441 0 0
0
0
4 VCO~
221 200 89 0 5 9
13 4 2 3 2 2
0
0 0 592 0
6 SQRVCO
20 -2 62 6
2 V1
35 -1 49 7
0
0
29 %D %%vd(%1,%2) %%vd(%3,%4) %M
0
13 alias:ASQRVCO
0
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
11 Signal Gen~
195 57 62 0 64 64
0 4 2 5 86 -10 10 9 0 0
0 0 0 0 0 0 0 1013276738 0 1036831949
990057071 1050253722 998445679 1065353216 1002740646 1069547520 1006834287 1056964608 1008981771 1075838976
1011129254 1082130432 1013276738 1036831949 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
20
0 0.014 0 0.1 0.002 0.3 0.004 1 0.006 1.5
0.008 0.5 0.01 2.5 0.012 4 0.014 0.1 0 0
0
0 0 848 0
4 0/4V
-15 -30 13 -22
2 V3
-7 -40 7 -32
0
0
77 %D %1 %2 DC 0 PWL( 0 100m 2m 300m 4m 1 6m 1.5 8m 500m 10m 2.5 12m 4 14m 100m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
7 Ground~
168 105 100 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
5 SAVE-
218 134 57 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
29 *Combine
*TRAN 0.000 10.00 5
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
7734 0 0
0
0
9 Resistor~
219 282 94 0 4 5
0 3 2 0 -1
0
0 0 880 270
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
6
1 3 3 0 0 8320 0 7 3 0 0 4
282 76
282 56
209 56
209 65
2 1 2 0 0 8192 0 4 5 0 0 3
88 67
105 67
105 94
1 0 2 0 0 0 0 1 0 0 5 2
193 151
193 134
4 0 2 0 0 0 0 3 0 0 5 2
209 119
209 134
2 2 2 0 0 8320 0 7 3 0 0 4
282 112
282 134
173 134
173 119
1 1 4 0 0 4224 0 4 3 0 0 3
88 57
173 57
173 65
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.014 5.6e-005 5.6e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
652 1079360 100 100 0 0
77 66 767 186
1 57 162 127
767 66
77 66
767 66
767 186
0 0
3e-005 0 5.4 0 3e-005 5.4
12385 0
4 1 0.05
0
668 8813120 100 100 0 0
77 66 767 186
0 319 800 572
767 66
77 66
767 66
767 186
0 0
0.014 0 5 -1 0.014 0.014
12409 0
4 2e-006 2
2
249 56
0 3 0 0 2	0 1 0 0
126 57
0 4 0 0 1	0 6 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
