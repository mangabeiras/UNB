CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 800 319
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\PROGRAM FILES\MICROCODE ENGINEERING\CIRCUITMAKER 6 PRO\BOM.DAT
0 7
0 66 800 319
12058624 0
1
6 Title:
5 Name:
0
0
0
11
3 PLL
219 236 101 0 8 17
0 7 8 8 2 3 5 6 4
3 PLL
0 0 15056 0
7 PLL100K
-29 8 20 16
4 PLL1
-40 -64 -12 -56
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
28 alias:XPLLX {Fc=100k Fr=50k}
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 -33686019
88 0 0 0 1 1 0 0
3 PLL
8953 0 0
0
0
2 +V
167 251 38 0 1 3
0 4
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 139 170 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 253 169 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
5 SAVE-
218 142 73 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
5 SAVE1
-11 -36 24 -28
0
0
11 *TRAN 0 5 0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
5394 0 0
0
0
11 Signal Gen~
195 35 70 0 64 64
0 7 2 3 86 -8 8 0 0 0
0 0 0 0 0 0 0 1203982336 1075838976 1075838976
1084227584 1176256512 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -33686019
20
0 100000 2.5 2.5 5 10000 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/5V
-14 -30 14 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SFFM(2.5 2.5 100k 5 10k)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
7 Ground~
168 85 169 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
10 Capacitor~
219 332 129 0 2 5
0 2 5
0
0 0 848 90
6 .002uF
12 0 54 8
2 C1
26 -10 40 -2
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
7 Ground~
168 332 172 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
9 Resistor~
219 253 133 0 3 5
0 2 3 -1
0
0 0 880 90
3 10k
7 0 28 8
2 R2
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 277 83 0 2 5
0 6 5
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
11
5 2 3 0 0 8320 0 1 10 0 0 3
241 101
253 101
253 115
8 1 4 0 0 8320 0 1 2 0 0 3
241 65
251 65
251 47
6 0 5 0 0 4224 0 1 0 0 5 2
241 92
332 92
7 1 6 0 0 4224 0 1 11 0 0 2
241 83
259 83
2 2 5 0 0 0 0 8 11 0 0 3
332 120
332 83
295 83
1 1 2 0 0 4096 0 8 9 0 0 2
332 138
332 166
1 1 7 0 0 4224 0 6 1 0 0 2
66 65
177 65
2 1 2 0 0 8320 0 6 7 0 0 3
66 75
85 75
85 163
3 2 8 0 0 4224 0 1 1 0 0 4
177 83
135 83
135 74
177 74
1 1 2 0 0 0 0 4 10 0 0 2
253 163
253 151
4 1 2 0 0 0 0 1 3 0 0 3
177 101
139 101
139 164
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.0002 2e-007 2e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
2 V1
0 10 1
0
0 0 0
5 -1 10 10 10 0 10 10 0
1508 1210432 100 100 0 0
0 0 0 0
0 66 161 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 2
0
1512 8550464 100 100 0 0
77 66 767 186
0 319 800 572
537 66
77 66
767 126
767 126
0 0
0.0002 0 0 0 0.0002 0.0002
13425 0
2 5e-005 5
4
154 65
0 7 0 -60 1	0 7 0 0
153 74
0 8 0 -31 3	0 9 0 0
245 83
0 6 0 1 1	0 4 0 0
244 101
0 3 0 39 1	0 1 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
