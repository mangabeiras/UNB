CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 300 100 3
0 66 520 452
7 5.000 V
7 5.000 V
3 GND
0 66 520 452
9961488 0
0
0
0
0
0
0
31
5 SAVE-
218 123 130 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
26 *Combine
*TRAN -250m 400m
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SAVE-
218 468 135 0 10 64
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
38 *Combine
*AC -1 550
*TRAN -250m 400m
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
10 Polar Cap~
219 271 270 0 2 64
0 5 4
10 Polar Cap~
0 0 336 0
6 3255pF
-19 12 23 20
2 C1
-7 5 7 13
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
10 Polar Cap~
219 356 270 0 2 64
0 4 6
10 Polar Cap~
0 0 336 0
6 1000pF
-21 12 21 20
2 C2
-8 4 6 12
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Capacitor~
219 452 135 0 2 64
0 6 7
10 Capacitor~
0 0 336 0
5 .47uF
-17 13 18 21
2 C3
-7 3 7 11
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
11 Signal Gen~
195 31 135 0 19 64
0 10 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1000593162
20
1 1000 0 0.005 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 16720 0
7 -5m/5mV
-24 -28 25 -20
2 V1
-7 -38 7 -30
0
0
37 %D %1 %2 DC 0 SIN(0 5m 1k 0 0) AC 1 0
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
7 Ground~
168 479 222 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
7 Ground~
168 372 203 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
7 Ground~
168 287 220 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
7 Ground~
168 239 220 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
7 Ground~
168 158 233 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
7 Ground~
168 111 233 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
7 Ground~
168 88 233 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
7 Ground~
168 72 163 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
2 +V
167 298 14 0 1 64
0 3
0
0 0 54128 0
5 +250V
11 8 46 16
6 Vplate
12 -4 54 4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
7 Triode~
219 169 130 0 3 64
0 9 10 5
7 Triode~
0 0 336 0
5 12AX7
13 17 48 25
2 Q1
26 6 40 14
0
0
14 %D %1 %2 %3 %S
0
0
0
7

0 1 2 3 1 2 3 -33686019
88 0 0 0 1 0 0 0
1 Q
4718 0 0
0
0
7 Triode~
219 298 133 0 3 64
0 11 13 12
7 Triode~
0 0 336 0
5 12AX7
13 -26 48 -18
2 Q2
30 2 44 10
0
0
14 %D %1 %2 %3 %S
0
0
0
7

0 1 2 3 1 2 3 -33686019
88 0 0 0 1 0 0 0
1 Q
3874 0 0
0
0
7 Triode~
219 383 92 0 3 64
0 3 11 8
7 Triode~
0 0 336 0
5 12AX7
15 -25 50 -17
2 Q3
30 1 44 9
0
0
14 %D %1 %2 %3 %S
0
0
0
7

0 1 2 3 1 2 3 -33686019
88 0 0 0 1 0 0 0
1 Q
6671 0 0
0
0
10 Capacitor~
219 88 197 0 2 64
0 10 2
10 Capacitor~
0 0 336 26894
4 36pF
-40 -3 -12 5
2 C4
19 -12 33 -4
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3789 0 0
0
0
10 Capacitor~
219 200 91 0 2 64
0 9 13
10 Capacitor~
0 0 336 0
4 .1uF
-15 -18 13 -10
2 C5
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
4871 0 0
0
0
10 Capacitor~
219 399 135 0 2 64
0 8 6
10 Capacitor~
0 0 336 0
5 .47uF
-17 13 18 21
2 C6
-7 3 7 11
0
0
11 %D %1 %2 %V
0
0
6 CAP0.2
5

0 1 2 1 2 -33686019
67 0 0 0 1 0 0 0
1 C
3750 0 0
0
0
9 Resistor~
219 269 248 0 2 64
0 5 4
9 Resistor~
0 0 368 0
5 1475k
-17 -12 18 -4
2 R1
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 354 248 0 2 64
0 4 6
9 Resistor~
0 0 368 0
3 75k
-10 -13 11 -5
2 R2
-7 -23 7 -15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 111 195 0 3 64
0 2 10 -1
9 Resistor~
0 0 368 90
5 47.5k
5 -2 40 6
2 R3
18 -12 32 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
9 Resistor~
219 158 193 0 3 64
0 2 5 -1
9 Resistor~
0 0 368 90
5 1.82k
9 0 44 8
2 R4
19 -12 33 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
9 Resistor~
219 239 186 0 3 64
0 2 13 -1
9 Resistor~
0 0 368 90
4 1Meg
6 -2 34 6
2 R5
13 -12 27 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
9 Resistor~
219 287 186 0 3 64
0 2 12 -1
9 Resistor~
0 0 368 90
2 1k
8 -2 22 6
2 R6
8 -12 22 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
5670 0 0
0
0
9 Resistor~
219 372 168 0 3 64
0 2 8 -1
9 Resistor~
0 0 368 90
4 100k
-38 -1 -10 7
2 R7
-31 -11 -17 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 169 62 0 4 64
0 9 3 0 1
9 Resistor~
0 0 368 90
4 300k
-34 -4 -6 4
2 R8
-27 -14 -13 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 298 66 0 4 64
0 11 3 0 1
9 Resistor~
0 0 368 90
4 100k
7 -4 35 4
2 R9
16 -9 30 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 479 179 0 3 64
0 2 7 -1
9 Resistor~
0 0 368 90
4 100k
-33 2 -5 10
3 R10
12 -13 33 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
33
1 0 3 0 0 8192 0 18 0 0 3 3
383 66
383 35
298 35
2 0 3 0 0 8320 0 29 0 0 3 3
169 44
169 35
298 35
1 2 3 0 0 0 0 15 30 0 0 2
298 23
298 48
0 0 4 0 0 4096 0 0 0 9 8 2
313 248
313 270
0 0 5 0 0 8320 0 0 0 28 7 4
158 165
214 165
214 260
241 260
0 0 6 0 0 4224 0 0 0 19 10 3
424 135
424 259
384 259
1 1 5 0 0 0 0 22 3 0 0 4
251 248
241 248
241 270
260 270
2 1 4 0 0 4224 0 3 4 0 0 2
277 270
345 270
1 2 4 0 0 0 0 23 22 0 0 2
336 248
287 248
2 2 6 0 0 0 0 23 4 0 0 4
372 248
384 248
384 270
362 270
2 2 7 0 0 8320 0 5 31 0 0 3
461 135
479 135
479 161
1 0 8 0 0 4096 0 21 0 0 21 2
390 135
372 135
1 0 9 0 0 4096 0 20 0 0 33 2
191 91
169 91
1 0 10 0 0 4096 0 19 0 0 30 2
88 188
88 130
2 1 2 0 0 4224 0 19 13 0 0 2
88 206
88 227
2 1 2 0 0 0 0 6 14 0 0 3
62 140
72 140
72 157
1 1 2 0 0 0 0 28 8 0 0 2
372 186
372 197
1 1 2 0 0 0 0 31 7 0 0 2
479 197
479 216
2 1 6 0 0 0 0 21 5 0 0 2
408 135
443 135
2 0 11 0 0 4224 0 18 0 0 32 2
357 92
298 92
2 3 8 0 0 4224 0 28 18 0 0 2
372 150
372 115
2 3 12 0 0 4224 0 27 17 0 0 2
287 168
287 156
2 0 13 0 0 4096 0 26 0 0 31 2
239 168
239 133
1 1 2 0 0 0 0 9 27 0 0 2
287 214
287 204
1 1 2 0 0 0 0 10 26 0 0 2
239 214
239 204
1 1 2 0 0 0 0 24 12 0 0 2
111 213
111 227
1 1 2 0 0 0 0 25 11 0 0 2
158 211
158 227
2 3 5 0 0 0 0 25 16 0 0 2
158 175
158 153
2 0 10 0 0 0 0 24 0 0 30 2
111 177
111 130
2 1 10 0 0 4224 0 16 6 0 0 2
143 130
62 130
2 2 13 0 0 8320 0 20 17 0 0 4
209 91
239 91
239 133
272 133
1 1 11 0 0 0 0 30 17 0 0 2
298 84
298 107
1 1 9 0 0 4224 0 29 16 0 0 2
169 80
169 104
1
-16 0 0 0 700 255 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
15 269 165 298
19 273 159 292
14 RIAA Amplifier
0
2073 0 1
0
0
6 Vplate
-10 300 2
0
0 0 0
10 2 10 20000
0 0.005 2e-005 2e-005 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
1936 1210432 100 100 0 0
77 66 287 126
0 66 140 136
287 66
77 66
287 66
287 126
0 0
0.00012 0.000100092 -7.7 -11.9 1.9908e-005 4.2
0 0
4 1 100
1
220 35
0 3 0 0 2	0 2 0 0
1916 8550464 100 100 0 0
77 66 287 126
320 66 640 259
287 66
77 66
287 66
287 126
0 0
0.005 0 0.8 -0.4 0.005 0.005
16 0
4 0.001 100
1
479 146
0 7 0 0 2	0 11 0 0
3464 4421696 100 100 0 0
98 66 294 126
320 259 640 452
258 66
98 66
294 66
294 66
0 0
19108.5 10 56 60.2 19098.5 19098.5
12387 0
4 5000 10000
1
479 150
0 7 0 0 2	0 11 0 0
0 0 100 100 0 0
77 66 293 126
0 0 0 0
293 66
77 66
293 66
293 126
0 0
1e+006 1 -3.55271e-015 -3.55271e-015 999999 999999
4211 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
