CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
10 70 30 70 9
0 66 640 259
8  5.000 V
8  5.000 V
3 GND
16666.7 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 259
9961482 0
0
0
0
0
0
0
53
5 SAVE-
218 55 159 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
5 SAVE1
-11 -36 24 -28
0
0
20 *TRAN -1.000 13.00 0
0
0
0
1

10 0
0 0 0 0 1 0 0 0
4 SAVE
8953 0 0
0
0
4 .IC~
207 115 188 0 1 3
0 5
0
0 0 53312 0
2 0V
-7 -15 7 -7
4 CMD1
-14 -25 14 -17
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
3 CMD
4441 0 0
0
0
2 +V
167 183 85 0 1 3
0 7
0
0 0 53600 0
3 +5V
12 -2 33 6
2 V1
15 -12 29 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
10 555 Timer~
219 125 150 0 8 17
0 2 5 3 8 6 5 4 7
10 555 Timer~
0 0 6464 0
3 555
-10 -23 11 -15
2 U2
-7 -33 7 -25
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 -33686019
88 0 0 0 1 1 0 0
1 U
6153 0 0
0
0
10 Polar Cap~
219 230 231 0 2 5
0 5 2
10 Polar Cap~
0 0 832 26894
4 .1uF
1 4 29 12
2 C1
10 -6 24 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
5394 0 0
0
0
10 Polar Cap~
219 177 230 0 2 5
0 6 2
10 Polar Cap~
0 0 832 26894
5 .01uF
7 4 42 12
2 C2
21 -6 35 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 0 0 0 1 1 0 0
1 C
7734 0 0
0
0
7 Ground~
168 129 267 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
4 4017
219 299 272 0 14 29
0 2 3 9 10 16 17 18 19 11
12 39 40 41 42
0
0 0 12512 0
4 4017
-14 -60 14 -52
2 U3
-7 -70 7 -62
0
15 DVDD=16;DGND=8;
102 %D [%16bi %8bi %1i %2i %3i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 13 14 15 3 2 4 7 10 1
5 6 9 11 12 13 14 15 3 2
4 7 10 1 5 6 9 11 12 -33686019
65 0 0 512 1 1 0 0
1 U
3747 0 0
0
0
9 3-In NOR~
219 415 385 0 4 21
0 11 16 10 13
0
0 0 96 0
4 4025
-14 -24 14 -16
3 U1C
-11 -34 10 -26
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 -33686019
65 0 0 0 3 3 2 0
1 U
3549 0 0
0
0
9 3-In NOR~
219 415 308 0 4 21
0 18 17 16 14
0
0 0 96 0
4 4025
-14 -24 14 -16
3 U1B
-11 -34 10 -26
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 -33686019
65 0 0 0 3 2 2 0
1 U
7931 0 0
0
0
9 3-In NOR~
219 417 230 0 4 21
0 11 19 18 15
0
0 0 96 0
4 4025
-14 -24 14 -16
3 U1A
-11 -34 10 -26
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 -33686019
65 0 0 0 3 1 2 0
1 U
9325 0 0
0
0
7 Ground~
168 797 402 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
13 Var Resistor~
219 668 338 0 3 7
0 7 24 24
13 Var Resistor~
0 0 320 0
7 500 40%
-25 8 24 16
2 R1
6 -22 20 -14
0
0
28 %DA %1 %2 200
%DB %2 %3 300
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 272 0 1 0 0 0
1 R
3834 0 0
0
0
4 LED~
171 764 388 0 2 5
10 25 2
0
0 0 96 90
4 LED2
10 -16 38 -8
2 D1
17 -26 31 -18
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3363 0 0
0
0
13 PNP Darling1~
219 735 365 0 3 7
0 25 22 23
13 PNP Darling1~
0 0 320 692
6 MPSA64
22 -5 64 3
2 Q1
27 -14 41 -6
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
88 0 242 256 1 1 0 0
1 Q
7668 0 0
0
0
10 Polar Cap~
219 624 366 0 2 5
0 7 22
10 Polar Cap~
0 0 320 270
5 100uF
10 -1 45 7
2 C3
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 -1 274 0 1 1 0 0
1 C
4718 0 0
0
0
7 Ground~
168 797 325 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3874 0 0
0
0
13 Var Resistor~
219 668 261 0 3 7
0 7 28 28
13 Var Resistor~
0 0 320 0
7 500 40%
-25 8 24 16
2 R2
6 -22 20 -14
0
0
28 %DA %1 %2 200
%DB %2 %3 300
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 272 0 1 0 0 0
1 R
6671 0 0
0
0
4 LED~
171 764 311 0 2 5
12 29 2
0
0 0 96 90
4 LED2
10 -16 38 -8
2 D2
17 -26 31 -18
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3789 0 0
0
0
13 PNP Darling1~
219 735 288 0 3 7
0 29 26 27
13 PNP Darling1~
0 0 320 692
6 MPSA64
22 -5 64 3
2 Q2
27 -14 41 -6
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
88 0 242 256 1 1 0 0
1 Q
4871 0 0
0
0
10 Polar Cap~
219 624 289 0 2 5
0 7 26
10 Polar Cap~
0 0 320 270
5 100uF
10 -1 45 7
2 C4
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 -1 274 0 1 1 0 0
1 C
3750 0 0
0
0
7 Ground~
168 795 174 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8778 0 0
0
0
7 Ground~
168 796 247 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
538 0 0
0
0
13 PNP Darling1~
219 735 134 0 3 7
0 33 32 34
13 PNP Darling1~
0 0 320 692
6 MPSA64
22 -5 64 3
2 Q3
27 -14 41 -6
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
88 0 242 256 1 1 0 0
1 Q
6843 0 0
0
0
13 Var Resistor~
219 669 106 0 3 7
0 7 30 30
13 Var Resistor~
0 0 320 0
7 500 40%
-25 8 24 16
2 R3
6 -22 20 -14
0
0
28 %DA %1 %2 200
%DB %2 %3 300
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 272 0 1 0 0 0
1 R
3136 0 0
0
0
4 LED~
171 763 159 0 2 5
21 33 2
0
0 0 96 90
4 LED3
10 -16 38 -8
2 D3
17 -26 31 -18
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5950 0 0
0
0
13 Var Resistor~
219 667 183 0 3 7
0 7 36 36
13 Var Resistor~
0 0 320 0
7 500 40%
-25 8 24 16
2 R4
6 -22 20 -14
0
0
28 %DA %1 %2 200
%DB %2 %3 300
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 272 0 1 0 0 0
1 R
5670 0 0
0
0
4 LED~
171 763 233 0 2 5
21 37 2
0
0 0 96 90
4 LED3
10 -16 38 -8
2 D4
17 -26 31 -18
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6828 0 0
0
0
13 PNP Darling1~
219 734 210 0 3 7
0 37 31 35
13 PNP Darling1~
0 0 320 692
6 MPSA64
22 -5 64 3
2 Q4
27 -14 41 -6
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
88 0 242 256 1 1 0 0
1 Q
6735 0 0
0
0
10 Polar Cap~
219 623 211 0 2 5
0 7 31
10 Polar Cap~
0 0 320 270
5 100uF
10 -1 45 7
2 C5
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 -1 274 0 1 1 0 0
1 C
8365 0 0
0
0
6 Diode~
219 480 385 0 2 5
0 20 13
6 Diode~
0 0 320 180
6 1N4148
-20 -18 22 -10
2 D5
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 -1 280 0 1 1 0 0
1 D
4132 0 0
0
0
6 Diode~
219 479 230 0 2 5
0 38 15
6 Diode~
0 0 320 180
6 1N4148
-20 -18 22 -10
2 D6
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 -1 280 0 1 1 0 0
1 D
4551 0 0
0
0
6 Diode~
219 479 308 0 2 5
0 21 14
6 Diode~
0 0 320 180
6 1N4148
-20 -18 22 -10
2 D7
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 -33686019
68 -1 280 0 1 1 0 0
1 D
3635 0 0
0
0
7 Ground~
168 243 321 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3973 0 0
0
0
10 Polar Cap~
219 349 145 0 2 5
0 7 9
10 Polar Cap~
0 0 320 270
5 .01uF
10 -1 45 7
2 C6
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 -1 274 0 1 1 0 0
1 C
3851 0 0
0
0
10 Polar Cap~
219 621 130 0 2 5
0 7 32
10 Polar Cap~
0 0 320 270
5 100uF
10 -1 45 7
2 C7
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 -33686019
67 -1 274 0 1 1 0 0
1 C
8383 0 0
0
0
9 Resistor~
219 31 201 0 3 5
0 2 3 -1
9 Resistor~
0 0 4960 90
3 10k
7 0 28 8
2 R5
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
9334 0 0
0
0
9 Resistor~
219 229 126 0 4 5
0 4 7 0 1
9 Resistor~
0 0 4960 90
3 250
7 0 28 8
2 R6
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 229 181 0 2 5
0 5 4
9 Resistor~
0 0 4960 90
3 250
4 -1 25 7
2 R7
8 -11 22 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3334 0 0
0
0
9 Resistor~
219 47 125 0 4 5
0 8 7 0 1
9 Resistor~
0 0 4960 90
2 2k
8 0 22 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 1 0 0
1 R
3559 0 0
0
0
9 Resistor~
219 715 338 0 2 5
0 24 23
9 Resistor~
0 0 352 0
2 47
-7 -12 7 -4
2 R9
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
984 0 0
0
0
9 Resistor~
219 582 363 0 3 5
0 7 22 1
9 Resistor~
0 0 352 270
3 47k
7 -5 28 3
3 R10
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
7557 0 0
0
0
9 Resistor~
219 531 385 0 2 5
0 20 22
9 Resistor~
0 0 352 0
3 47k
-11 -14 10 -6
3 R11
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
3146 0 0
0
0
9 Resistor~
219 715 261 0 2 5
0 28 27
9 Resistor~
0 0 352 0
2 47
-7 -12 7 -4
3 R12
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
5687 0 0
0
0
9 Resistor~
219 582 286 0 3 5
0 7 26 1
9 Resistor~
0 0 352 270
3 47k
7 -5 28 3
3 R13
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
7939 0 0
0
0
9 Resistor~
219 531 308 0 2 5
0 21 26
9 Resistor~
0 0 352 0
3 47k
-11 -14 10 -6
3 R14
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
3308 0 0
0
0
9 Resistor~
219 719 106 0 2 5
0 30 34
9 Resistor~
0 0 352 0
2 47
-7 -12 7 -4
3 R15
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
3408 0 0
0
0
9 Resistor~
219 714 183 0 2 5
0 36 35
9 Resistor~
0 0 352 0
2 47
-7 -12 7 -4
3 R16
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
9773 0 0
0
0
9 Resistor~
219 581 208 0 3 5
0 7 31 1
9 Resistor~
0 0 352 270
3 47k
7 -5 28 3
3 R17
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
691 0 0
0
0
9 Resistor~
219 580 128 0 3 5
0 7 32 1
9 Resistor~
0 0 352 270
3 47k
7 -5 28 3
3 R18
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
7834 0 0
0
0
9 Resistor~
219 531 151 0 2 5
0 38 32
9 Resistor~
0 0 352 0
3 47k
-11 -14 10 -6
3 R19
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
3588 0 0
0
0
9 Resistor~
219 530 230 0 2 5
0 38 31
9 Resistor~
0 0 352 0
3 47k
-11 -14 10 -6
3 R20
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
4528 0 0
0
0
9 Resistor~
219 348 199 0 2 5
0 9 12
9 Resistor~
0 0 352 270
4 1Meg
8 -5 36 3
3 R21
-10 -22 11 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 -1 271 0 1 1 0 0
1 R
3303 0 0
0
0
82
0 2 3 0 0 12416 0 0 8 11 0 4
31 167
10 167
10 299
267 299
2 0 4 0 0 4096 0 39 0 0 3 2
229 163
229 149
7 1 4 0 0 8320 0 4 38 0 0 4
157 150
157 149
229 149
229 144
1 0 5 0 0 4096 0 2 0 0 14 2
115 200
115 208
2 0 2 0 0 4096 0 6 0 0 12 2
176 237
176 250
1 5 6 0 0 4224 0 6 4 0 0 3
176 220
176 168
157 168
1 0 2 0 0 0 0 7 0 0 12 2
129 261
129 250
2 0 7 0 0 8192 0 40 0 0 17 3
47 107
47 106
183 106
4 1 8 0 0 4224 0 4 40 0 0 3
93 168
47 168
47 143
1 0 2 0 0 8192 0 37 0 0 12 3
31 219
31 228
68 228
3 2 3 0 0 0 0 4 37 0 0 3
93 159
31 159
31 183
1 2 2 0 0 12416 0 4 5 0 0 5
93 141
68 141
68 250
229 250
229 238
1 0 5 0 0 4096 0 5 0 0 15 2
229 221
229 208
2 0 5 0 0 12416 0 4 0 0 15 4
93 150
82 150
82 208
202 208
6 1 5 0 0 0 0 4 39 0 0 5
157 159
202 159
202 208
229 208
229 199
2 0 7 0 0 0 0 38 0 0 17 3
229 108
229 106
183 106
1 8 7 0 0 0 0 3 4 0 0 3
183 94
183 141
157 141
3 0 9 0 0 8320 0 8 0 0 33 4
267 317
256 317
256 165
348 165
1 1 2 0 0 0 0 8 34 0 0 3
261 290
243 290
243 315
4 3 10 0 0 8320 0 8 9 0 0 4
331 326
348 326
348 394
402 394
9 1 11 0 0 8320 0 8 9 0 0 4
331 281
368 281
368 376
402 376
10 2 12 0 0 8320 0 8 53 0 0 3
331 272
348 272
348 217
4 2 13 0 0 4224 0 9 31 0 0 2
454 385
470 385
4 2 14 0 0 4224 0 10 33 0 0 2
454 308
469 308
4 2 15 0 0 4224 0 11 32 0 0 2
456 230
469 230
3 0 16 0 0 4096 0 10 0 0 29 2
402 317
358 317
2 6 17 0 0 4224 0 10 8 0 0 2
403 308
331 308
1 7 18 0 0 4224 0 10 8 0 0 2
402 299
331 299
2 5 16 0 0 8320 0 9 8 0 0 4
403 385
358 385
358 317
331 317
3 0 18 0 0 0 0 11 0 0 28 3
404 239
388 239
388 299
2 8 19 0 0 8320 0 11 8 0 0 4
405 230
378 230
378 290
331 290
1 0 11 0 0 0 0 11 0 0 21 3
404 221
368 221
368 281
2 1 9 0 0 0 0 35 53 0 0 2
348 152
348 181
1 1 20 0 0 4224 0 43 31 0 0 2
513 385
490 385
1 1 21 0 0 4224 0 46 33 0 0 2
513 308
489 308
2 1 2 0 0 0 0 14 12 0 0 3
777 389
797 389
797 396
2 0 22 0 0 4096 0 16 0 0 39 2
623 373
623 385
2 0 22 0 0 0 0 42 0 0 39 2
582 381
582 385
2 2 22 0 0 4224 0 43 15 0 0 4
549 385
699 385
699 365
711 365
1 0 7 0 0 0 0 16 0 0 42 2
623 356
623 338
1 0 7 0 0 0 0 42 0 0 42 2
582 345
582 338
1 0 7 0 0 8192 0 13 0 0 71 3
650 338
562 338
562 106
2 3 23 0 0 4224 0 41 15 0 0 3
733 338
743 338
743 343
2 0 24 0 0 4224 0 13 0 0 45 3
666 326
690 326
690 338
3 1 24 0 0 0 0 13 41 0 0 2
686 338
697 338
1 1 25 0 0 8320 0 15 14 0 0 3
743 387
743 389
757 389
2 1 2 0 0 0 0 19 17 0 0 3
777 312
797 312
797 319
2 0 26 0 0 4096 0 21 0 0 50 2
623 296
623 308
2 0 26 0 0 0 0 45 0 0 50 2
582 304
582 308
2 2 26 0 0 4224 0 46 20 0 0 4
549 308
699 308
699 288
711 288
1 0 7 0 0 0 0 21 0 0 53 2
623 279
623 261
1 0 7 0 0 0 0 45 0 0 53 2
582 268
582 261
1 0 7 0 0 0 0 18 0 0 42 2
650 261
562 261
2 3 27 0 0 4224 0 44 20 0 0 3
733 261
743 261
743 266
2 0 28 0 0 4224 0 18 0 0 56 3
666 249
690 249
690 261
3 1 28 0 0 0 0 18 44 0 0 2
686 261
697 261
1 1 29 0 0 8320 0 20 19 0 0 3
743 310
743 312
757 312
2 1 2 0 0 0 0 28 23 0 0 3
776 234
796 234
796 241
2 1 2 0 0 0 0 26 22 0 0 3
776 160
795 160
795 168
1 0 7 0 0 0 0 35 0 0 71 2
348 135
348 106
1 0 7 0 0 0 0 50 0 0 71 2
580 110
580 106
1 0 7 0 0 0 0 36 0 0 71 2
620 120
620 106
2 0 30 0 0 4224 0 25 0 0 64 3
667 94
694 94
694 106
3 1 30 0 0 0 0 25 47 0 0 2
687 106
701 106
2 0 31 0 0 4096 0 30 0 0 67 2
622 218
622 230
2 0 31 0 0 0 0 49 0 0 67 2
581 226
581 230
2 2 31 0 0 4224 0 52 29 0 0 4
548 230
698 230
698 210
710 210
1 0 7 0 0 0 0 30 0 0 70 2
622 201
622 183
1 0 7 0 0 0 0 49 0 0 70 2
581 190
581 183
1 0 7 0 0 0 0 27 0 0 42 2
649 183
562 183
1 0 7 0 0 4224 0 25 0 0 16 2
651 106
229 106
2 0 32 0 0 4096 0 36 0 0 74 2
620 137
620 151
2 0 32 0 0 0 0 50 0 0 74 2
580 146
580 151
2 2 32 0 0 12416 0 24 51 0 0 4
711 134
697 134
697 151
549 151
1 1 33 0 0 8320 0 24 26 0 0 3
743 156
743 160
756 160
2 3 34 0 0 4224 0 47 24 0 0 3
737 106
743 106
743 112
2 3 35 0 0 4224 0 48 29 0 0 3
732 183
742 183
742 188
2 0 36 0 0 4224 0 27 0 0 79 3
665 171
689 171
689 183
3 1 36 0 0 0 0 27 48 0 0 2
685 183
696 183
1 1 37 0 0 8320 0 29 28 0 0 3
742 232
742 234
756 234
0 1 38 0 0 4224 0 0 51 82 0 3
505 230
505 151
513 151
1 1 38 0 0 0 0 32 52 0 0 2
489 230
512 230
1
-24 0 0 0 700 255 0 0 0 3 2 1 34
5 Arial
0 0 0 22
258 72 532 112
265 76 528 104
22 Multi-Chrome Projector
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.0003 6e-007 6e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2852 1210432 100 100 0 0
77 66 617 126
11 164 151 234
617 66
77 66
617 66
617 126
0 0
0 0 0 0 0 0
0 0
4 1 2
1
733 338
0 23 0 0 1	0 43 0 0
3480 8526400 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 86
617 96
0 0
0 0 0 0 0 0
13433 0
2 5e-005 5
4
187 299
0 3 0 21 3	0 1 0 0
506 385
0 20 0 0 1	0 34 0 0
504 308
0 21 0 -11 1	0 35 0 0
501 230
0 38 0 -30 1	0 82 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
