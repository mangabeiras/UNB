CircuitMaker Text
4
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 1e+012
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 100 0
0 66 640 236
0 236 640 452
159383552 0
0
0
0
0
0
0
9
5 SCOPE
12 593 22 0 4 
0 9 99 49 0 0
0 0 -7968 0
3 TP1
-11 -4 10 4
0
0
0
11 .PLOT V(%1)
0
2

0 1 0 
86 0 0 0 0 0 0 0
1 V
8953 0 0 0
5 SCOPE
12 553 22 0 4 
0 8 99 50 0 0
0 0 -7968 0
3 TP2
-11 -4 10 4
0
0
0
11 .PLOT V(%1)
0
2

0 1 0 
86 0 0 0 0 0 0 0
1 V
4441 0 0 0
5 SCOPE
12 514 22 0 5 
0 7 99 51 48 0 0
0 0 -7968 0
3 TP3
-11 -4 10 4
0
0
0
11 .PLOT V(%1)
0
2

0 1 0 
86 0 0 0 0 0 0 0
1 V
3618 0 0 0
5 SCOPE
12 475 22 0 5 
0 6 99 52 49 0 0
0 0 -7968 0
3 TP4
-11 -4 10 4
0
0
0
11 .PLOT V(%1)
0
2

0 1 0 
86 0 0 0 0 0 0 0
1 V
6153 0 0 0
5 SCOPE
12 436 23 0 5 
0 5 99 53 50 0 0
0 0 -7968 0
3 TP5
-11 -4 10 4
0
0
0
11 .PLOT V(%1)
0
2

0 1 0 
86 0 0 0 0 0 0 0
1 V
5394 0 0 0
5 SCOPE
12 395 23 0 5 
0 4 99 54 51 0 0
0 0 -7968 0
3 TP6
-11 -4 10 4
0
0
0
11 .PLOT V(%1)
0
2

0 1 0 
86 0 0 0 0 0 0 0
1 V
7734 0 0 0
5 SCOPE
12 353 23 0 5 
0 3 99 55 52 0 0
0 0 -7968 0
3 TP7
-11 -4 10 4
0
0
0
11 .PLOT V(%1)
0
2

0 1 0 
86 0 0 0 0 0 0 0
1 V
9914 0 0 0
5 SCOPE
12 210 28 0 5 
0 2 99 56 53 0 0
0 0 -7968 0
3 TP8
-11 -4 10 4
0
0
0
11 .PLOT V(%1)
0
2

0 1 0 
86 0 0 0 0 0 0 0
1 V
3747 0 0 0
10 Ascii Key~
169 271 39 0 12 
0 9 8 7 6 5 4 3 2 0 
0 116 0 0
0 0 20512 0
0
0
0
0
0
0
9

0 1 2 3 4 5 6 7 8 0 
0 0 0 0 0 0 0 0
0
3549 0 0 0
8
8 1 2 0 0 8320 0 9 8 0 0 4
250 63
250 77
210 77
210 40
7 1 3 0 0 8320 0 9 7 0 0 4
256 63
256 130
353 130
353 35
1 6 4 0 0 8320 0 6 9 0 0 4
395 35
395 121
262 121
262 63
5 1 5 0 0 8320 0 9 5 0 0 4
268 63
268 112
436 112
436 35
1 4 6 0 0 8320 0 4 9 0 0 4
475 34
475 105
274 105
274 63
3 1 7 0 0 8320 0 9 3 0 0 4
280 63
280 95
514 95
514 34
1 2 8 0 0 8320 0 2 9 0 0 4
553 34
553 85
286 85
286 63
1 1 9 0 0 8320 0 9 1 0 0 4
292 63
292 77
593 77
593 34
1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 133
6 9 206 133
10 13 202 109
133 Select the Key symbol 
by clicking on it. Run 
the simulation and 
type on the keyboard 
to display binary data 
waveforms.
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
