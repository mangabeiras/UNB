CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 3
0 66 444 342
7 5.000 V
7 5.000 V
3 GND
0 66 444 342
-1031798782 0
2
0
0
0
0
0
13
13 Logic Switch~
5 151 99 0 2 3
169 13 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 S1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 151 118 0 2 3
192 12 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 S2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 151 158 0 2 3
0 10 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 S3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 150 177 0 2 3
0 9 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 S4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 151 198 0 2 3
0 8 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 S5
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 151 218 0 2 3
0 7 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 S6
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 231 58 0 2 3
0 15 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 S7
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 230 78 0 2 3
0 14 -99
0
0 0 20592 0
2 0V
-7 -16 7 -8
2 S8
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
7 Ground~
168 50 199 0 1 3
0 16
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
3549 0 0
0
0
9 Data Seq~
170 48 105 0 17 21
0 17 18 19 20 21 22 23 11 24
25 13 1 20 1 1 0 33
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -54 10 -46
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
0
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
7931 0 0
0
0
AAAAABAAABAAABAAABAAABAAABAAABAAABAAABAAABAAAAAAAAAAAAAAAAAAAAAAAA
12 Hex Display~
7 384 43 0 4 9
10 2 3 4 5
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -52 17 -44
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9325 0 0
0
0
14 Logic Display~
6 325 64 0 1 3
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
7 74LS168
8 223 159 0 14 29
0 13 12 11 10 9 8 7 14 15
6 5 4 3 2
0
0 0 12528 0
8 74LS168A
-28 -60 28 -52
2 U1
-7 -70 7 -62
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 -33686019
65 0 0 0 1 1 0 0
1 U
3834 0 0
0
0
14
1 14 2 0 0 8320 0 11 13 0 0 3
393 67
393 195
255 195
2 13 3 0 0 8320 0 11 13 0 0 3
387 67
387 186
255 186
3 12 4 0 0 8320 0 11 13 0 0 3
381 67
381 177
255 177
4 11 5 0 0 8320 0 11 13 0 0 3
375 67
375 168
255 168
1 10 6 0 0 4224 0 12 13 0 0 3
325 82
325 159
261 159
1 7 7 0 0 8320 0 6 13 0 0 4
163 218
179 218
179 195
191 195
1 6 8 0 0 12416 0 5 13 0 0 4
163 198
170 198
170 186
191 186
1 5 9 0 0 4224 0 4 13 0 0 2
162 177
191 177
1 4 10 0 0 4224 0 3 13 0 0 4
163 158
180 158
180 168
191 168
8 3 11 0 0 4224 0 10 13 0 0 2
80 141
191 141
1 2 12 0 0 8320 0 2 13 0 0 3
163 118
163 132
185 132
1 1 13 0 0 8320 0 1 13 0 0 4
163 99
175 99
175 123
185 123
1 8 14 0 0 8320 0 8 13 0 0 4
242 78
269 78
269 123
261 123
1 9 15 0 0 8320 0 7 13 0 0 4
243 58
285 58
285 132
255 132
6
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 12
93 171 135 214
97 175 136 210
12 Preset
Data
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 15
300 12 356 51
304 16 357 51
15 Terminal
Count
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 7
154 47 214 69
158 51 226 71
7 Up/Down
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 5
27 150 68 173
31 154 69 174
5 Clock
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 14
84 90 139 128
88 94 140 129
14 Count
Enables
-13 0 0 0 400 0 0 0 0 3 2 1 18
15 Times New Roman
0 0 0 13
139 66 221 89
143 70 222 90
13 Parallel Load
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 2e-005 8e-008 8e-008 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 100 100 0 0
77 66 617 126
0 0 0 0
617 66
77 66
617 66
617 126
0 0
0.0008333 0 0.6 -0.6 0.0008333 0.0008333
16 0
0 0.0002 10
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
0.0005 0 1.2 -1.2 0.0005 2.4
16 0
0 5e-006 10
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
2000 1 2.38857 0 1999 1999
16 0
0 500 1000
0
0 0 100 100 0 0
98 66 296 126
0 0 0 0
296 66
98 66
296 66
296 126
0 0
1e+006 1 -3.55271e-015 0 999999 999999
12403 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
